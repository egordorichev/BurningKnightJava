 3 M         Z                                                                            %                                                                                                                   &                                                                                              '                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       !                                                                                                                                                                                                                                                                                                     !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 !                                                                                                                                              #                                                                         +                                                                 +                                                                 +                                                                 +                                                                 *                                                                         )                                                  )                                                                                *                                                                       *                                                                       *                                                                       )                                                                                                                         "                                                                        �        �       �       �        �       �                 "                                                                                 �        �        �        �        �       �                 #                                                                         �        �                         �        �                 #                                                                         �       �                        �       �                 #                                                                     �        �        �        �        �        �                         "                                                                      �       �       �       �       �        �                #                                                                                                    '                                                                +                                                                        )                                                                               *                                                                         *                                                                 '                                                 &                                                                                                                %                                                                                                         %                                                                                                                 &                                                                                                         %                                                                                                                 &                                                                                                               %                                                                                                             %                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             &                                                                                            oM o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . R o l l i n g S p i k e R o o m     , N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . L i n e E n t r a n c e R o o m  <  F  F o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s h o p . Q u a d S h o p R o o m  =  D J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . H a l f R o o m C h a s m  2  < H o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s p e c i a l . N p c S a v e R o o m  ? ( K J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . G o l d S e c r e t R o o m  % # ,H o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . b o s s . S i m p l e B o s s R o o m   %  T o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . t r e a s u r e . C o r n e r l e s s T r e a s u r e R o o m %  1  K o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . F i l l e d R o m b R o o m  <  H N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . B o s s E n t r a n c e R o o m 	 F  J S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . E m p t y C o n n e c t i o n R o o m  ,  2 O o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . C h a s m T u n n e l R o o m      S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . C h a s m C o n n e c t i o n R o o m  : " ? J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . T u n n e l R o o m %  (    
  	
 
	

 
    N e n t i t y . t r a p . R o l l i n g S p i k e  z   A�       e n t i t y . t r a p . R o l l i n g S p i k e  T  P��       e n t i t y . t r a p . R o l l i n g S p i k e  �  �A�       e n t i t y . l e v e l . e n t i t i e s . E n t r a n c e   �  
  e n t i t y . l e v e l . e n t i t i e s . S l a b   1  � e n t i t y . i t e m . I t e m H o l d e r   3  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b       e n t i t y . l e v e l . e n t i t i e s . S l a b   a  � e n t i t y . i t e m . I t e m H o l d e r   f  �E o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . p e t . o r b i t a l . N a n o O r b i t a l       e n t i t y . l e v e l . e n t i t i e s . S l a b   1   e n t i t y . i t e m . I t e m H o l d e r   3  #F o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . w e a p o n . s w o r d . M o r n i n g S t a r        e n t i t y . l e v e l . e n t i t i e s . S l a b   a   e n t i t y . i t e m . I t e m H o l d e r   c  #P o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . a c c e s s o r y . e q u i p p a b l e . D e f e n s e E m b l e m   
    " e n t i t y . c r e a t u r e . n p c . B l u e S h o p k e e p e r   `  0 ( (        e n t i t y . i t e m . I t e m H o l d e r   d  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r   $  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . l e v e l . e n t i t i e s . D o o r        6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C " B e n t i t y . c r e a t u r e . n p c . T r a d e r     P 
 
        d e n t i t y . i t e m . I t e m H o l d e r    `2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �  `2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �  p2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r    �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �  `2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d       ' e n t i t y . l e v e l . e n t i t i e s . c h e s t . W o o d e n C h e s t  �   ` @ o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . w e a p o n . s p e a r . S p e a r          e n t i t y . l e v e l . e n t i t i e s . P o r t a l   �  x  e n t i t y . c r e a t u r e . f x . F i r e f l y   �   e n t i t y . c r e a t u r e . f x . F i r e f l y   �  � e n t i t y . c r e a t u r e . f x . F i r e f l y   �  N e n t i t y . c r e a t u r e . f x . F i r e f l y   7  " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  @  �  e n t i t y . c r e a t u r e . f x . F i r e f l y  �   v e n t i t y . c r e a t u r e . f x . F i r e f l y  t   Z e n t i t y . c r e a t u r e . f x . F i r e f l y  �   �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `   0" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b      0" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `   �  e n t i t y . c r e a t u r e . f x . F i r e f l y  m  K e n t i t y . c r e a t u r e . f x . F i r e f l y  b  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  p" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  p   � e n t i t y . c r e a t u r e . f x . F i r e f l y  p   � e n t i t y . l e v e l . e n t i t i e s . D o o r  p  �      , e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �        e n t i t y . l e v e l . e n t i t i e s . D o o r   �  �      < e n t i t y . l e v e l . e n t i t i e s . D o o r          B e n t i t y . l e v e l . e n t i t i e s . D o o r   �  0  6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C  C e n t i t y . l e v e l . e n t i t i e s . D o o r   �  X   < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . B u r n i n g K e y 
 F e n t i t y . l e v e l . e n t i t i e s . D o o r  �        2 e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �     ; e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �      ? e n t i t y . l e v e l . e n t i t i e s . D o o r  T   �    %  e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �       e n t i t y . l e v e l . e n t i t i e s . D o o r  p   �     '  e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  �  �         e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �  ` 
 
        e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  P  ` 
 
       % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  �  0         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �  � 
 
        e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �   � 
 
        e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  �   0         e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  �   �        e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  @  +         e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  ^  9  
      % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  _  �         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  `  @ 
 
        e n t i t y . i t e m . I t e m H o l d e r  �  �O o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . c o n s u m a b l e . s c r o l l . S c r o l l O f U p g r a d e        e n t i t y . i t e m . I t e m H o l d e r  ?  L2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . i t e m . I t e m H o l d e r  3  o< o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . e n t i t i e s . C o i n        e n t i t y . i t e m . I t e m H o l d e r  b  �6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C       