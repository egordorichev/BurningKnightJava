   	 s e t t i n g s _ f u l l s c r e e n f a l s e s e t t i n g s _ g o r e t r u e s e t t i n g s _ q u a l i t y 1 s e t t i n g s _ v s y n c t r u e s e t t i n g s _ s f x 0 . 5 s e t t i n g s _ m u s i c 0 . 5 s e t t i n g s _ u i s f x t r u e s e t t i n g s _ b l o o d t r u e s e t t i n g s _ s c r e e n s h a k e 0 . 7