 � >                                                           ~                                                                        }                                                                       R                                                                                                                                                                                                    P                                                                                                                                                                                                                                                                                               P                                                                                                                                                                                                                                                                                           P                                                                                                                                                                                                                                                                                                                                                   O                                                                                                                                                                                                                                                                                                                                                                                                                  O                                                                                                                                                                                                                                                                                                                                                                                            P                                                                                                                                                                                                                                                                                                                                  X                                                                                                                                                                                                                                                                                                                                                           X                                                                                                                                                                                                                                                                                                                     W                                                                                                                                                                                                                                                                                                      V                                                                                                                                                                                                                                                                                                                                 	                                                                                                      0                                                                                                                                                                                                                                                                                                                                                              	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    
                                                                                                                                                                                                 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �        �       �       �       �        �                                                                                                                         !                                                                                                                                                                                                                                                                                                                                                                                                                                        �       �       �       �        �        �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             	�       �        �       �        �        �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     
�       �       �       �        �       �                                                           (                                                                                                                                                                                                                                                                                                                                                                                                                                                                       	        �        �       �       �        �        �                2                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       	�        �        �       �       �        �                         1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
�       �       �        �       �        �                         1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          C                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    C                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 A                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          C                                                                                                                                                                                                                                                                                                                                                                                                                                                               C                                                                                                                                                                                                                                                                                                                                                                                                                              C                                                                                                                                                                                                                                                                                 \                                                                                                                                                                                              	                                                                               [                                                                                                                                                                                                                                                                                             \                                                                                                                                                                                        	                                                                             Z                                                                                                                                                                                                                                                                                            [                                                                                                                                                                                                                                                                                                [                                                                                                                                                                                        	                                                                                [                                                                                                                                                                                             
                                                                           Y                                                                                                                                                                                                                                                      Z                                                                                                                                                                                                                     \                                                                                                                                                                                                                                                  ]                                                                                                                                                    �                                      �                 �                                          �                        ~                                                                                                                                                                                                                                                                }                                                                                                                                                   ~                                                                                                                         ~                                                                                                          hM o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . D o u b l e C o r n e r R o o m "  , * D o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . P a d R o o m k  }  G o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . C i r c l e R o o m Y  g  N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . S m a l l A d d i t i o n R o o m O  Y  J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . C a v y C h a s m R o o m 0  E " J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . b o s s . C o l l u m n s B o s s R o o m    . J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . E n t r a n c e R o o m }  � 	  S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . t r e a s u r e . B r o k e L i n e T r e a s u r e R o o m $ 2 , < D o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . B o m b R o o m O  V R o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . R i n g C o n n e c t i o n R o o m g  k  R o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . R i n g C o n n e c t i o n R o o m J  O  P o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . S p i k e d T u n n e l R o o m E  J  P o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . S p i k e d T u n n e l R o o m ,  0 ! S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . E m p t y C o n n e c t i o n R o o m   "   R o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . R i n g C o n n e c t i o n R o o m * * / 2    		
		


      D e n t i t y . l e v e l . e n t i t i e s . E n t r a n c e     J ' e n t i t y . l e v e l . e n t i t i e s . c h e s t . W o o d e n C h e s t  �  p M o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . a c c e s s o r y . e q u i p p a b l e . P o i s o n R i n g        e n t i t y . i t e m . I t e m H o l d e r  3  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . i t e m . I t e m H o l d e r  3  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . i t e m . I t e m H o l d e r  3  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . c r e a t u r e . f x . F i r e f l y  D  a e n t i t y . c r e a t u r e . f x . F i r e f l y  }  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  0  @" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  P  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �   � e n t i t y . c r e a t u r e . f x . F i r e f l y  |  " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �   P" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  p  0  e n t i t y . c r e a t u r e . f x . F i r e f l y  r  � e n t i t y . c r e a t u r e . f x . F i r e f l y    � e n t i t y . c r e a t u r e . f x . F i r e f l y  K  � e n t i t y . c r e a t u r e . f x . F i r e f l y    x" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �    e n t i t y . c r e a t u r e . f x . F i r e f l y  �  0 e n t i t y . c r e a t u r e . f x . F i r e f l y  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b    �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  � e n t i t y . l e v e l . e n t i t i e s . D o o r  $  �     "   e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �      + *  e n t i t y . l e v e l . e n t i t i e s . D o o r  �        ,    e n t i t y . l e v e l . e n t i t i e s . D o o r  �   �     }   e n t i t y . l e v e l . e n t i t i e s . D o o r  �   �     k   e n t i t y . l e v e l . e n t i t i e s . D o o r  �   p     Y   e n t i t y . l e v e l . e n t i t i e s . D o o r  t   `     g   e n t i t y . l e v e l . e n t i t i e s . D o o r  �       O   e n t i t y . l e v e l . e n t i t i e s . D o o r  T  @     E   e n t i t y . l e v e l . e n t i t i e s . D o o r    �     0   e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �       e n t i t y . l e v e l . e n t i t i e s . D o o r  �        + 2  e n t i t y . l e v e l . e n t i t i e s . D o o r  �       J    e n t i t y . c r e a t u r e . m o b . d e s e r t . M u m m y  p  � 
 
       $ e n t i t y . c r e a t u r e . m o b . c o m m o n . M o v i n g F l y  �  �         $ e n t i t y . c r e a t u r e . m o b . c o m m o n . M o v i n g F l y  `  �         $ e n t i t y . c r e a t u r e . m o b . c o m m o n . M o v i n g F l y  p  �         $ e n t i t y . c r e a t u r e . m o b . c o m m o n . M o v i n g F l y  0  �         # e n t i t y . c r e a t u r e . m o b . D i a g o n a l S h o t F l y  4  @         # e n t i t y . c r e a t u r e . m o b . d e s e r t . S k e l e t o n  �  @         $ e n t i t y . c r e a t u r e . m o b . c o m m o n . M o v i n g F l y     `         ' e n t i t y . c r e a t u r e . m o b . d e s e r t . A r c h e o l o g i s t  �    
 
       $ e n t i t y . c r e a t u r e . m o b . c o m m o n . M o v i n g F l y  �   �         $ e n t i t y . c r e a t u r e . m o b . c o m m o n . M o v i n g F l y  �   �         $ e n t i t y . c r e a t u r e . m o b . c o m m o n . M o v i n g F l y  P   �         $ e n t i t y . c r e a t u r e . m o b . c o m m o n . M o v i n g F l y  @   �         ' e n t i t y . c r e a t u r e . m o b . d e s e r t . A r c h e o l o g i s t    P 
 
       ' e n t i t y . c r e a t u r e . m o b . d e s e r t . A r c h e o l o g i s t  0   
 
        e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  0   �         $ e n t i t y . c r e a t u r e . m o b . c o m m o n . M o v i n g F l y  p   �         $ e n t i t y . c r e a t u r e . m o b . c o m m o n . M o v i n g F l y  0   �         $ e n t i t y . c r e a t u r e . m o b . c o m m o n . M o v i n g F l y             $ e n t i t y . c r e a t u r e . m o b . c o m m o n . M o v i n g F l y  `            & e n t i t y . c r e a t u r e . m o b . c o m m o n . D i a g o n a l F l y  �   �         # e n t i t y . c r e a t u r e . m o b . d e s e r t . S k e l e t o n      �         ' e n t i t y . c r e a t u r e . m o b . d e s e r t . A r c h e o l o g i s t    0 
 
       # e n t i t y . c r e a t u r e . m o b . D i a g o n a l S h o t F l y  )  q         & e n t i t y . c r e a t u r e . m o b . c o m m o n . D i a g o n a l F l y    �         # e n t i t y . c r e a t u r e . m o b . D i a g o n a l S h o t F l y    �         ' e n t i t y . c r e a t u r e . m o b . d e s e r t . A r c h e o l o g i s t  �    
 
        e n t i t y . i t e m . I t e m H o l d e r  o   �< o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . e n t i t i e s . C o i n       