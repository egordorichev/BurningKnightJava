    s e t t i n g s _ g o r e t r u e s e t t i n g s _ q u a l i t y 1 U N L O C K _ D E W _ V I A L t r u e h i d e _ m i n i m a p t r u e s e t t i n g s _ b l t r u e s e t t i n g s _ v s y n c t r u e
 l a s t _ c l a s s 0 s e t t i n g s _ u i s f x t r u e s e t t i n g s _ b l o o d t r u e s e t t i n g s _ s a 8 s e t t i n g s _ f u l l s c r e e n f a l s e n u m _ f i r e _ o u t 1 D I E _ A C H I E V E M E N T t r u e s e t t i n g s _ c u r s o r c u r s o r - s m a l l R E A C H _ D E S E R T _ A C H I E V E M E N T t r u e s e t t i n g s _ s m t r u e s e t t i n g s _ r o t a t e _ c u r s o r f a l s e f i n i s h e d _ t u t o r i a l t r u e s e t t i n g s _ s f x 0 . 7 5 s e t t i n g s _ s t t r u e s e t t i n g s _ m u s i c 0 . 5 d e a t h s 1 s e t t i n g s _ s c r e e n s h a k e 0 . 7 T U T O R I A L _ D O N E _ A C H I E V E M E N T t r u e