 6 J         8                                                  .                                                                         ,                                                                                  ,                                                                         .                                                                                                           (                                                                                                                                         &                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                #                                                                                                                                                   !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        $                                                                                                                                     �       �        �        �        �        �        �                                                                                                                                            �        �       �        �       �        �        �                                                                                                                            �        �       �        �        �       �        �                         #                                                         �        �        �       �        �        �        �                %                                                 �        �       �       �       �        �       �                         $                                                         �        �       �        �       �        �       �                 #                                                                                                                            "                                                                                                                                                                     "                                                                                                                                                                   !                                                                                                                                                           "                                                                                                                                                                 !                                                                                                                                                                                                                                                                                                                                                           "                                                                                                                                                                 !                                                                                                                                                                                 !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �        �        �        �        �        �        �                .�       �        �        �        �        �        �                 -        �        �        �        �       �        �        �                 .�        �        �        �       �       �        �                        -�        �       �       �        �       �       �                 .�        �        �        �       �        �        �                .                                  �P o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . C i r c l e E n t r a n c e R o o m      R o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . V e r t i c a l S p i k e T r a p R o o m   & 4 0 Q o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . t r e a s u r e . C o l l u m n T r e a s u r e R o o m   	  H o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . b o s s . S i m p l e B o s s R o o m  0 4 A K o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . M i x e d S e c r e t R o o m  A ! HJ o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . G o l d S e c r e t R o o m ,  4 &E o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . R o m b R o o m 
    I o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . T r i a n g l e R o o m   , " N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . B o s s E n t r a n c e R o o m     S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . E m p t y C o n n e c t i o n R o o m # " ) & O o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . C h a s m T u n n e l R o o m     O o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . C h a s m T u n n e l R o o m 	       
 	 
 	 		
 


   I e n t i t y . l e v e l . e n t i t i e s . E n t r a n c e  �   �  e n t i t y . t r a p . R o l l i n g S p i k e  !  ��   ��  ! e n t i t y . l e v e l . e n t i t i e s . c h e s t . M i m i c   P   `           e n t i t y . i t e m . I t e m H o l d e r  �  `2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . i t e m . I t e m H o l d e r  �   2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . i t e m . I t e m H o l d e r  �  P2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . i t e m . I t e m H o l d e r  �   6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C        e n t i t y . i t e m . I t e m H o l d e r  �  @6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C        e n t i t y . i t e m . I t e m H o l d e r  �  02 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �  P2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . c r e a t u r e . f x . H e a r t F x  �  0 e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  P 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  0 
 
       e n t i t y . i t e m . I t e m H o l d e r  �   2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  3   2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  3  02 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r     2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �  02 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �   2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �  P2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �  2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . l e v e l . e n t i t i e s . P o r t a l  �   � " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �   � e n t i t y . c r e a t u r e . f x . F i r e f l y  3  � e n t i t y . c r e a t u r e . f x . F i r e f l y   _   Y e n t i t y . c r e a t u r e . f x . F i r e f l y   E   � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  1 e n t i t y . c r e a t u r e . f x . F i r e f l y  V  A e n t i t y . c r e a t u r e . f x . F i r e f l y  �  ;" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  0  " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �    " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  0    e n t i t y . c r e a t u r e . f x . F i r e f l y  ,  - e n t i t y . c r e a t u r e . f x . F i r e f l y  �  2 e n t i t y . c r e a t u r e . f x . F i r e f l y    $" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  0 e n t i t y . c r e a t u r e . f x . F i r e f l y      e n t i t y . c r e a t u r e . f x . F i r e f l y    p e n t i t y . c r e a t u r e . f x . F i r e f l y  g  � e n t i t y . c r e a t u r e . f x . F i r e f l y  h  " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �   �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �   " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �   e n t i t y . c r e a t u r e . f x . F i r e f l y  �   �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �   � e n t i t y . c r e a t u r e . f x . F i r e f l y  h  H e n t i t y . c r e a t u r e . f x . F i r e f l y  `  @" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  @  P  e n t i t y . c r e a t u r e . f x . F i r e f l y  Z   �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b      e n t i t y . l e v e l . e n t i t i e s . D o o r  �          e n t i t y . l e v e l . e n t i t i e s . D o o r  �   �       e n t i t y . l e v e l . e n t i t i e s . D o o r  �   �   < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . B u r n i n g K e y   e n t i t y . l e v e l . e n t i t i e s . D o o r  p  X      ' & e n t i t y . l e v e l . e n t i t i e s . D o o r    �      1 0 e n t i t y . l e v e l . e n t i t i e s . D o o r   �   p     	  e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �       e n t i t y . l e v e l . e n t i t i e s . D o o r  �        ( " e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f    � 
 
        e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  p  � 
 
        e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  0  p 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  �  �         e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n   �  �        % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t   �  �         e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n             e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  @            e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �    
 
        e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �   � 
 
        e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n     �         e n t i t y . i t e m . I t e m H o l d e r  !  �O o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . c o n s u m a b l e . s c r o l l . S c r o l l O f U p g r a d e        e n t i t y . i t e m . I t e m H o l d e r   �  >< o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . e n t i t i e s . C o i n       