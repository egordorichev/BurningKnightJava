 * <         U                                                                                                                                                                                                                                                                                                                                                                                                                                                                 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           �     �     �     �     �     �      �                                                                                                                                                                                                                                                          �     �      �      �      �      �      �      �                                                                                                                                                                                                                                                            �      �            �     �     �             �                                                                                                                                                                                                                                                            �            �                                                                                                                                                                    �     �             �                                                                                                                                                                                                                                                                                   �      �      �                                                                                                                                                                                                                       �      �      �                                                                                                                                                                                                           �                                                                                               �     �      �                                                                                                                                                                                                                                                           �      �     �                                                                                                                     �      �                          �     �      �      �                                                                                                             �     �     �                                                                                                                   �      �                    �      �      �      �     �                                                                                                                                                                                                                                                       �      �      �      �     �     �     �      �      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           �     �     �                                                                                                                                                                                                                                                                                               �      �     �                                                                                                                                                                                                                                                                                            �     �      �     �                                                                                                                                                                                                                                                                                             �      �     �      �                                                                                                                                                                                                                                                                                               �            �                                                                                                                                                                                                                                                                                             �            �                                                                                                                                                                                                                                                                                �     �     �      �     �                                                                                                                                                                                                                                                                          �             �     �     �      �                                                                                                                                                                                                                                                                �      �       �                                                                                                                                                                                                                                                                                          �       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               
                                                                                                                                                                                                                < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m  &  3 < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m  	   < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m   &  < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m   '  < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m    & < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m  3  9     % e n t i t y . l e v e l . e n t i t i e s . D o o r   �  X      
 & e n t i t y . l e v e l . e n t i t i e s . D o o r   �  X        e n t i t y . l e v e l . e n t i t i e s . D o o r   �  (       3' e n t i t y . l e v e l . e n t i t i e s . c h e s t . W o o d e n C h e s t  �   �  e n t i t y . c r e a t u r e . p l a y e r . S p a w n     h   ' 9 e n t i t y . l e v e l . e n t i t i e s . T r e e  �   L e n t i t y . l e v e l . e n t i t i e s . T r e e  0   � e n t i t y . l e v e l . e n t i t i e s . T r e e  @   | e n t i t y . l e v e l . e n t i t i e s . S t o n e  �  l
 p r o p _ s t o n e  e n t i t y . l e v e l . e n t i t i e s . S t o n e     L
 p r o p _ s t o n e  e n t i t y . l e v e l . e n t i t i e s . S t o n e   �   � p r o p _ b i g _ s t o n e e n t i t y . l e v e l . e n t i t i e s . S t o n e  @   <
 p r o p _ s t o n e e n t i t y . l e v e l . e n t i t i e s . T r e e  0   , e n t i t y . l e v e l . e n t i t i e s . T r e e   `   e n t i t y . l e v e l . e n t i t i e s . S t o n e  �   � p r o p _ b i g _ s t o n e e n t i t y . l e v e l . e n t i t i e s . T r e e  �   \ e n t i t y . l e v e l . e n t i t i e s . T r e e   �  � e n t i t y . l e v e l . e n t i t i e s . T r e e   �   e n t i t y . l e v e l . e n t i t i e s . S t o n e   0  l p r o p _ h i g h _ s t o n e e n t i t y . l e v e l . e n t i t i e s . S t o n e  �   �
 p r o p _ s t o n e  e n t i t y . l e v e l . e n t i t i e s . S t o n e      �
 p r o p _ s t o n e! e n t i t y . l e v e l . e n t i t i e s . R o l l T r i g g e r  �  ' e n t i t y . l e v e l . e n t i t i e s . c h e s t . W o o d e n C h e s t   �  � M o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . c o n s u m a b l e . p o t i o n . H e a l i n g P o t i o n        ' e n t i t y . l e v e l . e n t i t i e s . c h e s t . W o o d e n C h e s t  @  , A o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . w e a p o n . g u n . R e v o l v e r             ! e n t i t y . l e v e l . e n t i t i e s . T u t o r i a l E n d   �  � e n t i t y . c r e a t u r e . f x . F i r e f l y    � e n t i t y . c r e a t u r e . f x . F i r e f l y   �  G e n t i t y . c r e a t u r e . f x . F i r e f l y     � e n t i t y . c r e a t u r e . f x . F i r e f l y   �   e n t i t y . c r e a t u r e . f x . F i r e f l y   U  - e n t i t y . c r e a t u r e . f x . F i r e f l y     l e n t i t y . c r e a t u r e . f x . F i r e f l y  D   � e n t i t y . c r e a t u r e . f x . F i r e f l y   �   e n t i t y . c r e a t u r e . f x . F i r e f l y   �   e n t i t y . c r e a t u r e . f x . F i r e f l y   �   e n t i t y . c r e a t u r e . f x . F i r e f l y   �  ; e n t i t y . c r e a t u r e . f x . H e a r t F x    �