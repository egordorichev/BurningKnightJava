    e n t i t y . c r e a t u r e . p l a y e r . P l a y e r  e  �        A o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . w e a p o n . g u n . R e v o l v e r              N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . a c c e s s o r y . e q u i p p a b l e . P o i s o n B o m b s      M o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . a c c e s s o r y . e q u i p p a b l e . B l a c k H e a r t    
   L o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . a c c e s s o r y . e q u i p p a b l e . B i g B u l l e t      L o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . a c c e s s o r y . e q u i p p a b l e . O l d M a n u a l                       A�       & e n t i t y . c r e a t u r e . m o b . b o s s . B u r n i n g K n i g h t����     2 2          