   ( s e t t i n g s _ g o r e t r u e U N L O C K _ B L A C K _ H E A R T t r u e U N L O C K _ D E W _ V I A L t r u e h i d e _ m i n i m a p f a l s e U N L O C K _ M I M I C _ T O T E M t r u e U N L O C K _ M E E T B O Y _ A X E t r u e F I N D _ M I M I C _ A C H I E V E M E N T t r u e	 n u m _ c o i n s 4 R E A C H _ D E S E R T _ A C H I E V E M E N T t r u e s e t t i n g s _ r o t a t e _ c u r s o r t r u e f i n i s h e d _ t u t o r i a l t r u e s e t t i n g s _ f f 0 . 5 s e t t i n g s _ m u s i c 0 . 5
 s e t t i n g s _ v f a l s e U N L O C K _ S A L E t r u e s e t t i n g s _ s c r e e n s h a k e 0 . 3 U N L O C K _ D I A M O N D t r u e s e t t i n g s _ f r f 0 . 5 n u m _ b u l l e t s _ r e f l e c t e d 2 s e t t i n g s _ q u a l i t y 2 s e t t i n g s _ b l f a l s e s e t t i n g s _ v s y n c t r u e
 l a s t _ c l a s s 0 s e t t i n g s _ s f f a l s e s e t t i n g s _ u i s f x t r u e U N L O C K _ M E E T B O Y t r u e s e t t i n g s _ b l o o d t r u e s e t t i n g s _ s a 0 s e t t i n g s _ f u l l s c r e e n f a l s e n u m _ f i r e _ o u t 1 s e t t i n g s _ c u r s o r c u r s o r - s t a n d a r t s e t t i n g s _ s m f a l s e n p c _ d _ s a v e d t r u e s e t t i n g s _ s f x 0 . 7 5 s e t t i n g s _ s t f a l s e E Q U I P _ A C C E S S O R Y _ A C H I E V E M E N T t r u e U N L O C K _ M I M I C _ S U M M O N E R t r u e s e t t i n g s _ c b 0 . 0 T U T O R I A L _ D O N E _ A C H I E V E M E N T t r u e n u m _ k e y s _ u s e d 0