_L     x                           V                                                      1                                                                                  0                                                                          1                                                                                                5                                                                                   ?                                                                                                /                                                                                                                                                                                                                                                                                                                                             	                                                                                                                                                                                                                                                  	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       
                                                                                                                                                                                                            /                                                                                                                                                  /                                                                                                                          
                                   *                                                                                                                                                                (                                                                                                                                                       (                                                                                                                                  (                                                                                                                                   '                                                                                                                                   '                                                                                                                                        (                                                                                          ,                                                                                               ,                                                                                                   ,                                                                                                                                               %                                                                                                                                                                    !�   �    �    �   �    �    �   �    �                                                                                                                                                   !    �    �   �    �   �   �    �    �    �                                                                                                                                                    !    �    �    �    �    �    �   �    �    �                                                                                                                                                     !    �   �    �    �    �   �    �   �    �                                                                                                                                                    !�    �   �    �    �    �   �    �    �                                                                                                                                                 "�   �    �    �    �    �    �    �    �                                                                                                                                                       !�    �    �    �   �    �    �    �   �                                                                                                                                              
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �    �    �    �    �    �   �                                                                                                                                                                              �    �    �    �   �    �   �                                                                                                                                                                                �    �    �    �    �    �    �                                                                                                                                                                                                                           �   �    �       �    �   �                                                                                                                                                                                         �    �    �    �    �   �    �   �   �    �    �                                         �   �    �   �   �   �    �                                                                                                                                                                  �    �   �    �   �    �    �    �    �    �    �                                        �    �    �   �    �    �    �                                                                                                                                                                                 �   �   �   �    �    �    �    �   �   �   �                                    �   �    �    �   �    �   �                	                                                                                                                                                                    �    �    �   �    �    �    �   �    �   �    �                                                       	                                                                                                                                                     	�    �    �    �    �    �    �    �    �   �    �                                                                                                 	                                                                                                                                                                 �    �    �   �    �    �    �    �   �    �   �                                                                                                
                                                                                	                                                                                                        �    �    �    �    �    �    �   �   �    �    �                                                                                               
                                                                                         
         �   �   �   �    �   �   �    �    �    �    �                                                                                                                                                                     '                                                                                                     	                                                                                  ,                                                                                                                                                                  ,                                                                                              	                                                                        +                                                                                                 	                                                                    ,                                                                                                                                                               ,                                                                                                                                                                                 *                                                                                                                         	                                                          +                                                                                                                   	                                                          ,                                                                                                                            	   	                                                 +                                                                                                                                                             ,                                                                                                                                        G                                                                                          I                                                                                 L                                                                       L                                                                M                                                                    V                               �N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . B o s s E n t r a n c e R o o m   #  E o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . H e a r t R o o m  "  *I o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . C o l l u m n s R o o m    + J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . E n t r a n c e R o o m , > 1 I  N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . t r e a s u r e . M a z e T r e a s u r e R o o m 8  H  G o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . P r i s o n R o o m D ) ] 8 N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . M i s s i n g C o r n e r R o o m 1 / ; > J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . G o l d S e c r e t R o o m  - " 5G o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . T u r r e t R o o m ; + D > H o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . b o s s . S i m p l e B o s s R o o m  	   K o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . i t e m . B r o k e L i n e I t e m R o o m 4  > + Q o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . t r e a s u r e . C o l l u m n T r e a s u r e R o o m  ! # - J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . C a v y C h a s m R o o m !  8  F o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s h o p . G o l d S h o p R o o m  1  :E o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . C a v e R o o m  5 ' D P o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . S p i k e d T u n n e l R o o m ' B , F S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . E m p t y C o n n e c t i o n R o o m  1  5 S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . E m p t y C o n n e c t i o n R o o m  +  1 J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . T u n n e l R o o m   ! 	 S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . C h a s m C o n n e c t i o n R o o m /  6  J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . T u n n e l R o o m > > E C E o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . C a v e R o o m 1 > > J 8 		
			 

	
   � e n t i t y . l e v e l . e n t i t i e s . E x i t     H  e n t i t y . c r e a t u r e . f x . H e a r t F x   C  p  e n t i t y . c r e a t u r e . f x . H e a r t F x   s  � e n t i t y . c r e a t u r e . f x . H e a r t F x   s  @ e n t i t y . c r e a t u r e . f x . H e a r t F x   3  0  e n t i t y . l e v e l . e n t i t i e s . E n t r a n c e  �  : ! e n t i t y . l e v e l . e n t i t i e s . c h e s t . M i m i c      �           e n t i t y . i t e m . I t e m H o l d e r  �  02 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �  02 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �   2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . t r a p . T u r r e t  �  �>��      e n t i t y . t r a p . T u r r e t  �   >��       e n t i t y . t r a p . T u r r e t  �  0>��       e n t i t y . t r a p . T u r r e t  �  `>��      e n t i t y . t r a p . T u r r e t  �  �>��      e n t i t y . t r a p . T u r r e t  �  �>��      e n t i t y . l e v e l . e n t i t i e s . S l a b  �   e n t i t y . i t e m . I t e m H o l d e r  �  O o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . c o n s u m a b l e . s c r o l l . S c r o l l O f U p g r a d e       % e n t i t y . l e v e l . e n t i t i e s . c h e s t . I r o n C h e s t  �  p M o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . a c c e s s o r y . e q u i p p a b l e . R e d B a l l o o n        e n t i t y . i t e m . I t e m H o l d e r   �  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r   �  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r   �  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . l e v e l . e n t i t i e s . S l a b   r  8 e n t i t y . i t e m . I t e m H o l d e r   t  ?2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b   
   e n t i t y . l e v e l . e n t i t i e s . S l a b   �  8 e n t i t y . i t e m . I t e m H o l d e r   �  ?6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C   
   e n t i t y . l e v e l . e n t i t i e s . S l a b   �  8 e n t i t y . i t e m . I t e m H o l d e r   �  BE o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . w e a p o n . s w o r d . L i g h t s a b e r   
     e n t i t y . l e v e l . e n t i t i e s . S l a b   �  8 e n t i t y . i t e m . I t e m H o l d e r   �  ?Q o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . a c c e s s o r y . e q u i p p a b l e . G r a v i t y B o o s t e r       e n t i t y . l e v e l . e n t i t i e s . S l a b   �  8 e n t i t y . i t e m . I t e m H o l d e r   �  =L o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . a c c e s s o r y . e q u i p p a b l e . F i r e B o o t s       e n t i t y . l e v e l . e n t i t i e s . S l a b    8 e n t i t y . i t e m . I t e m H o l d e r    <R o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . a c c e s s o r y . e q u i p p a b l e . P e n e t r a t i o n R u n e   
  $ e n t i t y . c r e a t u r e . n p c . O r a n g e S h o p k e e p e r   p  p        " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �  e n t i t y . c r e a t u r e . f x . F i r e f l y  (  F e n t i t y . c r e a t u r e . f x . F i r e f l y  �   e n t i t y . c r e a t u r e . f x . F i r e f l y  �  f" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �   0" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  p   0" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  0 " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `  � " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  P  0" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  0" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  @  @" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  `" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     p" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �   " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     �  e n t i t y . c r e a t u r e . f x . F i r e f l y  �   e n t i t y . c r e a t u r e . f x . F i r e f l y  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b   �   �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �   �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b   �  � " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  b   e n t i t y . c r e a t u r e . f x . F i r e f l y  t  :" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  P  �  e n t i t y . c r e a t u r e . f x . F i r e f l y  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �  e n t i t y . c r e a t u r e . f x . F i r e f l y  E   � e n t i t y . c r e a t u r e . f x . F i r e f l y  �   � e n t i t y . c r e a t u r e . f x . F i r e f l y   �  G e n t i t y . c r e a t u r e . f x . F i r e f l y   �  A e n t i t y . c r e a t u r e . f x . F i r e f l y   �  2 e n t i t y . c r e a t u r e . f x . F i r e f l y  .  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  `" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `   " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �   �  e n t i t y . c r e a t u r e . f x . F i r e f l y  ;  @" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �    e n t i t y . c r e a t u r e . f x . F i r e f l y  U  1 e n t i t y . c r e a t u r e . f x . F i r e f l y  �  G" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  `" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `  � " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �  e n t i t y . l e v e l . e n t i t i e s . D o o r  �         	    e n t i t y . l e v e l . e n t i t i e s . D o o r  p  �         + e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �        * e n t i t y . l e v e l . e n t i t i e s . D o o r   �  �      	    e n t i t y . l e v e l . e n t i t i e s . D o o r    �       1 ? e n t i t y . l e v e l . e n t i t i e s . D o o r  �  @       , D e n t i t y . l e v e l . e n t i t i e s . D o o r  �   �       8  e n t i t y . l e v e l . e n t i t i e s . D o o r  D          D 0 e n t i t y . l e v e l . e n t i t i e s . D o o r  P  �        5 > e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �      
  < + e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �        ? > e n t i t y . l e v e l . e n t i t i e s . D o o r  �   �     	    	 e n t i t y . l e v e l . e n t i t i e s . D o o r  P  h     
   5  e n t i t y . l e v e l . e n t i t i e s . D o o r  @   �        4  e n t i t y . l e v e l . e n t i t i e s . D o o r     �       !  e n t i t y . l e v e l . e n t i t i e s . D o o r  @  H         5 e n t i t y . l e v e l . e n t i t i e s . D o o r  t  0       ' C e n t i t y . l e v e l . e n t i t i e s . D o o r  �         > A& e n t i t y . c r e a t u r e . m o b . h a l l . F r e e z i n g C l o w n  �  P         e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n   �           % e n t i t y . c r e a t u r e . m o b . h a l l . B u r n i n g C l o w n  @  0         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �  �          e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f   �           % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t    :        ' e n t i t y . c r e a t u r e . m o b . h a l l . S t a b b i n g K n i g h t  @           e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �  p          e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  P             e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  @  @         " e n t i t y . c r e a t u r e . m o b . h a l l . B o s s T h i e f  @  @         # e n t i t y . c r e a t u r e . m o b . h a l l . I n v i s T h i e f  �           % e n t i t y . c r e a t u r e . m o b . h a l l . B u r n i n g C l o w n     �         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f     �         ' e n t i t y . c r e a t u r e . m o b . h a l l . S t a b b i n g K n i g h t  0            e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  @           & e n t i t y . c r e a t u r e . m o b . h a l l . F r e e z i n g C l o w n  P            e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  `  �          e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  �  �        ' e n t i t y . c r e a t u r e . m o b . h a l l . S t a b b i n g K n i g h t  �  0         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f     P         # e n t i t y . c r e a t u r e . m o b . h a l l . I n v i s T h i e f  �  p          e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t      
 
      % e n t i t y . c r e a t u r e . m o b . h a l l . B u r n i n g C l o w n  �  `         e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  �  P        e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �  �          e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  `            e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  b  { 
 
      ' e n t i t y . c r e a t u r e . m o b . h a l l . S t a b b i n g K n i g h t  p  �        ' e n t i t y . c r e a t u r e . m o b . h a l l . S t a b b i n g K n i g h t  �  �        % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  �  `         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �  �         ' e n t i t y . c r e a t u r e . m o b . h a l l . S t a b b i n g K n i g h t     �         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f     �          e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f      �       
  e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  �   �        & e n t i t y . c r e a t u r e . m o b . h a l l . F r e e z i n g C l o w n  0   �         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �   �       	  e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  P   �         e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  p   � 
 
      & e n t i t y . c r e a t u r e . m o b . h a l l . F r e e z i n g C l o w n  �   �        ' e n t i t y . c r e a t u r e . m o b . h a l l . S t a b b i n g K n i g h t     �        % e n t i t y . c r e a t u r e . m o b . h a l l . B u r n i n g C l o w n  �  �         e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  0  �         e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �   
 
      # e n t i t y . c r e a t u r e . m o b . h a l l . I n v i s T h i e f  0  �         e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  p           e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  P           % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  w  k        % e n t i t y . c r e a t u r e . m o b . h a l l . B u r n i n g C l o w n  �          # e n t i t y . c r e a t u r e . m o b . h a l l . I n v i s T h i e f               e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  0  @        % e n t i t y . c r e a t u r e . m o b . h a l l . B u r n i n g C l o w n  0  p        e n t i t y . i t e m . I t e m H o l d e r  �  c< o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . e n t i t i e s . C o i n       