 � /         �                                                                                                                                                                                o                                                                                                                                                                                                                                                          h                                                                                                                                                                                                                                                                                                 b                                                                                                                                                                                                                                                                                                                                                                      3                                                                                                                                                                                                                                                                                                                                                                                                                                                                     2                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   1                                                                                                       #                                                                                                                                                                                                                                                                                                                                                                                                                                          8                                                                                     "                                                                                                                                                                                                                                                                                                                                                                                                                                                                  5                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            
                                                                                                                                                                                                                                                 (                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                +                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           
                                                                                                                                              0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           1                                                                                                                                                                                                                                    
                                                                                                                                                                                                                                                                                                                                                                                                                 1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                2                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           L                                                                                                                                                                                                                                                                                                                                                                                                                                                                                j                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     j                                                                                                                                                                                                                                                                                                                                                                                                                                                             h                                                                                                                                                                                                                                                                                                                                                                                                                 i                                                                                                                                                                                                                                                                                                                                                                                  j                                                                                                                                                                                                                                                                                                                                                                                          h                                                                                                                                                                                                                                                                                                                                                                                                                                      j                                                                                                                                                                                                                                                                                                                                                                                                                                          i                                                                                                                                                                                                                                                                                                                                                                                                                                          i                                                                                                                                                            
                                                                                                                                                                                                                                                        i                                                                                                                                                                                              	                                                                                                                                                                                                                                                   i                                                                                                                                                                                               
                                                                                                                                                                                                                                               i                                                                                                                                                                                                                                                                                                                                                                                                          t                                                                                                                                                                                                                                                                                                                            t                                                                                            
                                                                                                                                                                                                                                                t                                                                                                    
                                                                                                                                                                                                                                                t                                                                                                                                                                                                                                                                                  �                                                                                                                                                                                                                                        �                                                                                                                                                                                                                                              �                                                                                                                                                                                                                                             �                                                                                                    [F o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . T u t o r i a l C h a s m R o o m      P o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . C i r c l e E n t r a n c e R o o m 	     J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . b o s s . C o l l u m n s B o s s R o o m �  � - H o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s p e c i a l . N p c S a v e R o o m s   ) G o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . C o r n e r R o o m '  1  F o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . C r o s s R o o m 1  G  E o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . R o m b R o o m S 	 a  K o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . C e n t e r W a l l R o o m h  s % G o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . C i r c l e R o o m y  �  T o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . t r e a s u r e . C o r n e r l e s s T r e a s u r e R o o m     K o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . M i x e d S e c r e t R o o m   	  U o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . B i g R i n g C o n n e c t i o n R o o m    '  R o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . R i n g C o n n e c t i o n R o o m G  K  S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . C h a s m C o n n e c t i o n R o o m K  S  J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . T u n n e l R o o m a  h  O o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . C h a s m T u n n e l R o o m s  y  U o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . B i g R i n g C o n n e c t i o n R o o m s  y  &   	 
	 
    Z e n t i t y . l e v e l . e n t i t i e s . E n t r a n c e   �   �  e n t i t y . l e v e l . e n t i t i e s . D o o r  �     6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C y "  e n t i t y . c r e a t u r e . n p c . T r a d e r  �  @ 
 
         d e n t i t y . c r e a t u r e . f x . H e a r t F x   3   @ e n t i t y . c r e a t u r e . f x . H e a r t F x   c   � e n t i t y . c r e a t u r e . f x . F i r e f l y   �   � e n t i t y . c r e a t u r e . f x . F i r e f l y   �   � e n t i t y . c r e a t u r e . f x . F i r e f l y   �   � e n t i t y . c r e a t u r e . f x . F i r e f l y   �   � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  � " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  p  0 e n t i t y . c r e a t u r e . f x . F i r e f l y  �   � e n t i t y . c r e a t u r e . f x . F i r e f l y  �   �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �    " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `   �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  0   � " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  P   �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  P  0 " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     @" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  `  e n t i t y . c r e a t u r e . f x . F i r e f l y  �  ) e n t i t y . c r e a t u r e . f x . F i r e f l y  �   � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  J" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �   �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �   � " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �   �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `   �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `   " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  0 " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  @  e n t i t y . c r e a t u r e . f x . F i r e f l y  m   �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b      P" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  P   `" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  0 " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  P " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y   i   q e n t i t y . c r e a t u r e . f x . F i r e f l y  [   � e n t i t y . c r e a t u r e . f x . F i r e f l y     � e n t i t y . c r e a t u r e . f x . F i r e f l y  D  " e n t i t y . c r e a t u r e . f x . F i r e f l y  z  6 e n t i t y . c r e a t u r e . f x . F i r e f l y  `  � e n t i t y . l e v e l . e n t i t i e s . D o o r     �        e n t i t y . l e v e l . e n t i t i e s . D o o r   �   �     
  e n t i t y . l e v e l . e n t i t i e s . D o o r  �   �        e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �    �  e n t i t y . l e v e l . e n t i t i e s . D o o r  `  �     v   e n t i t y . l e v e l . e n t i t i e s . D o o r  t   �    '   e n t i t y . l e v e l . e n t i t i e s . D o o r     �    1   e n t i t y . l e v e l . e n t i t i e s . D o o r  t   �    G   e n t i t y . l e v e l . e n t i t i e s . D o o r         a   e n t i t y . l e v e l . e n t i t i e s . D o o r  4       S   e n t i t y . l e v e l . e n t i t i e s . D o o r  4  �    s   e n t i t y . l e v e l . e n t i t i e s . D o o r  �       h   e n t i t y . l e v e l . e n t i t i e s . D o o r  4  0    s   e n t i t y . l e v e l . e n t i t i e s . D o o r  �  0    y   e n t i t y . l e v e l . e n t i t i e s . D o o r  �   �    K  % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  �   �         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  @   �         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �   �        & e n t i t y . c r e a t u r e . m o b . c o m m o n . D i a g o n a l F l y  e   x         e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  �     	 	      $ e n t i t y . c r e a t u r e . m o b . c o m m o n . M o v i n g F l y  �  P        % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t      �         e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �   �         e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  �  @ 	 	      " e n t i t y . c r e a t u r e . m o b . c o m m o n . C o i n M a n  �   �        & e n t i t y . c r e a t u r e . m o b . c o m m o n . D i a g o n a l F l y  �  @         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f      �         e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  �   � 	 	       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t      
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t    0 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f    p 2 2       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �           e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t      � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �   �         e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t     p         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f             % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  p           e n t i t y . i t e m . I t e m H o l d e r  �  �6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C        e n t i t y . c r e a t u r e . f x . H e a r t F x  �   �' e n t i t y . l e v e l . e n t i t i e s . c h e s t . W o o d e n C h e s t  p  0  e n t i t y . i t e m . I t e m H o l d e r        2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r        2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r        2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r        2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r        2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �   �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d       