 2 V         e                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       �             �                                                                                                                                                                                                                                                                                                                     �             �      �     �                                                                                                                                                                                                                                                                                                                    �      �      �      �      �                                                                                                                                                                                                                                                                                                                  �                    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �            �                                                                                                                                                                                                                                                                                                                                         �      �      �      �                                                                                                                                                                                                                                                                                                                  �      �      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �< o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m 
 D  O < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m 
 8  D < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m  #  8 < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m    # < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m   . # < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m   .      ' e n t i t y . l e v e l . e n t i t i e s . D o o r  T  �      % ' e n t i t y . l e v e l . e n t i t i e s . c h e s t . W o o d e n C h e s t  �  H  e n t i t y . c r e a t u r e . p l a y e r . S p a w n  �   � e n t i t y . l e v e l . e n t i t i e s . T r e e  p   � e n t i t y . l e v e l . e n t i t i e s . T r e e  �   ` e n t i t y . l e v e l . e n t i t i e s . T r e e  @   � e n t i t y . l e v e l . e n t i t i e s . T r e e  �   � e n t i t y . l e v e l . e n t i t i e s . T r e e       e n t i t y . l e v e l . e n t i t i e s . T r e e      � e n t i t y . l e v e l . e n t i t i e s . T r e e  �   � e n t i t y . l e v e l . e n t i t i e s . T r e e  P   � e n t i t y . l e v e l . e n t i t i e s . T r e e  `    e n t i t y . l e v e l . e n t i t i e s . T r e e  �    e n t i t y . l e v e l . e n t i t i e s . T r e e  �    e n t i t y . l e v e l . e n t i t i e s . T r e e     ` e n t i t y . l e v e l . e n t i t i e s . T r e e  0  p e n t i t y . l e v e l . e n t i t i e s . T r e e     � e n t i t y . l e v e l . e n t i t i e s . T r e e  �  ` e n t i t y . l e v e l . e n t i t i e s . S t o n e     P
 p r o p _ s t o n e e n t i t y . l e v e l . e n t i t i e s . S t o n e   `  �
 p r o p _ s t o n e  e n t i t y . l e v e l . e n t i t i e s . S t o n e     
 p r o p _ s t o n e  e n t i t y . l e v e l . e n t i t i e s . S t o n e  �  @
 p r o p _ s t o n e  e n t i t y . l e v e l . e n t i t i e s . S t o n e  �  0
 p r o p _ s t o n e  e n t i t y . l e v e l . e n t i t i e s . S t o n e      � p r o p _ h i g h _ s t o n e e n t i t y . l e v e l . e n t i t i e s . S t o n e     p p r o p _ h i g h _ s t o n e e n t i t y . l e v e l . e n t i t i e s . S t o n e  @   � p r o p _ h i g h _ s t o n e e n t i t y . l e v e l . e n t i t i e s . S t o n e  �   � p r o p _ h i g h _ s t o n e e n t i t y . l e v e l . e n t i t i e s . S t o n e      � p r o p _ b i g _ s t o n e e n t i t y . l e v e l . e n t i t i e s . S t o n e  @  P p r o p _ b i g _ s t o n e e n t i t y . l e v e l . e n t i t i e s . S t o n e  P  � p r o p _ b i g _ s t o n e  e n t i t y . c r e a t u r e . f x . F i r e f l y   �  � e n t i t y . c r e a t u r e . f x . F i r e f l y   �  h e n t i t y . c r e a t u r e . f x . F i r e f l y  S  1 e n t i t y . c r e a t u r e . f x . F i r e f l y  !  � e n t i t y . c r e a t u r e . f x . F i r e f l y    � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y     e n t i t y . c r e a t u r e . f x . F i r e f l y  �   � e n t i t y . c r e a t u r e . f x . H e a r t F x   �  �