    e n t i t y . c r e a t u r e . p l a y e r . P l a y e r  �          F o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . w e a p o n . s w o r d . M o r n i n g S t a r        M o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . c o n s u m a b l e . p o t i o n . H e a l i n g P o t i o n                         A�     & e n t i t y . c r e a t u r e . m o b . b o s s . B u r n i n g K n i g h t         d d         