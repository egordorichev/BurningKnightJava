 [ 2         �                         W�        �        �        �        �       �                 T�        �        �        �        �        �                 T�       �        �        �       �        �                         R        �        �        �        �        �        �                        S�       �       �        �       �        �                T�        �       �       �        �       �                        S�        �        �       �        �       �                 T�        �        �        �        �       �                 T�        �        �        �       �       �                 S                                                           U                                                     P                                                                                 P                                                                          P                                                                   P                                                                                                                                                                             2                                                                                                                                                                                                                                                                            *                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �        �        �        �        �        �        �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �       �        �        �        �        �        �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �        �       �       �        �       �        �                                                                                                                                                                                                                                                                                                                                                                                                     �        �        �        �        �        �       �                                                                                                                                                                                                                                                                                                                                                                                      �        �        �        �        �       �       �                                                                                                                                                                                                                       �        �        �        �        �        �        �                                                                                                                                                                     /�       �        �        �       �        �       �                                                                                                                                                     0�       �        �        �        �        �        �                                                                                                                                                             /�        �       �       �       �        �        �                                                                                                                                                   5                                                                                                                                                     J                                                                                                                                     J                                                                                                                                             I                                                                                                                                               H                                                                                                                                                J                                                                                                                                       J                                                                                                              �E o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . H e a r t R o o m B  J )G o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . C i r c l e R o o m 4  B $ E o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . H e a r t R o o m D  K M o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . R o l l i n g S p i k e R o o m    0 N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . L i n e E n t r a n c e R o o m N  U   H o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . b o s s . S i m p l e B o s s R o o m   , % S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . t r e a s u r e . B r o k e L i n e T r e a s u r e R o o m     N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . B o s s E n t r a n c e R o o m U  Y  F o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . C r o s s R o o m E  N  U o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . B i g R i n g C o n n e c t i o n R o o m =  E  J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . T u n n e l R o o m ,  4 " S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . C h a s m C o n n e c t i o n R o o m    " S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . E m p t y C o n n e c t i o n R o o m       	
 
	 		

   J e n t i t y . c r e a t u r e . f x . H e a r t F x  3    e n t i t y . c r e a t u r e . f x . H e a r t F x  �   e n t i t y . c r e a t u r e . f x . H e a r t F x  S     e n t i t y . c r e a t u r e . f x . H e a r t F x  S    e n t i t y . c r e a t u r e . f x . H e a r t F x  3    e n t i t y . c r e a t u r e . f x . H e a r t F x  �   �  e n t i t y . c r e a t u r e . f x . H e a r t F x  �   � e n t i t y . c r e a t u r e . f x . H e a r t F x  �   @  e n t i t y . t r a p . R o l l i n g S p i k e   �  ���  �    e n t i t y . t r a p . R o l l i n g S p i k e   k   A�  �    e n t i t y . t r a p . R o l l i n g S p i k e   �  0��  �    e n t i t y . t r a p . R o l l i n g S p i k e   k  `A�  �    e n t i t y . t r a p . R o l l i n g S p i k e   �  ���  �    e n t i t y . t r a p . R o l l i n g S p i k e   k  �A�  �    e n t i t y . l e v e l . e n t i t i e s . E n t r a n c e  !  Z ' e n t i t y . l e v e l . e n t i t i e s . c h e s t . G o l d e n C h e s t   �  ` @ o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . w e a p o n . g u n . C h o p p e r             e n t i t y . l e v e l . e n t i t i e s . P o r t a l  p    e n t i t y . c r e a t u r e . f x . F i r e f l y  A  A e n t i t y . c r e a t u r e . f x . F i r e f l y  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  P  � " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b    � e n t i t y . c r e a t u r e . f x . F i r e f l y  z   | e n t i t y . c r e a t u r e . f x . F i r e f l y  l   E e n t i t y . c r e a t u r e . f x . F i r e f l y    � e n t i t y . c r e a t u r e . f x . F i r e f l y  ;  | e n t i t y . c r e a t u r e . f x . F i r e f l y    w e n t i t y . c r e a t u r e . f x . F i r e f l y  �  v" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  @ " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b    �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `   e n t i t y . c r e a t u r e . f x . F i r e f l y  �  ;" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `  P  e n t i t y . c r e a t u r e . f x . F i r e f l y  ,  ^ e n t i t y . c r e a t u r e . f x . F i r e f l y    W e n t i t y . c r e a t u r e . f x . F i r e f l y    F e n t i t y . c r e a t u r e . f x . F i r e f l y    G" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  @  ` e n t i t y . c r e a t u r e . f x . F i r e f l y    � e n t i t y . c r e a t u r e . f x . F i r e f l y    �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  � " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     � " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  0  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `   e n t i t y . c r e a t u r e . f x . F i r e f l y  @  � e n t i t y . c r e a t u r e . f x . F i r e f l y  V  � e n t i t y . c r e a t u r e . f x . F i r e f l y  K  � e n t i t y . c r e a t u r e . f x . F i r e f l y  W  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `  � e n t i t y . l e v e l . e n t i t i e s . D o o r  D  �     4  e n t i t y . l e v e l . e n t i t i e s . D o o r    h      A  e n t i t y . l e v e l . e n t i t i e s . D o o r  $  �       e n t i t y . l e v e l . e n t i t i e s . D o o r  T    < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . B u r n i n g K e y U  e n t i t y . l e v e l . e n t i t i e s . D o o r  �  P     N  e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �     ,  e n t i t y . l e v e l . e n t i t i e s . D o o r  t        ! e n t i t y . l e v e l . e n t i t i e s . D o o r  t  �       e n t i t y . l e v e l . e n t i t i e s . D o o r  $  �       e n t i t y . l e v e l . e n t i t i e s . D o o r  T  P     E & e n t i t y . c r e a t u r e . m o b . c o m m o n . D i a g o n a l F l y    �        & e n t i t y . c r e a t u r e . m o b . c o m m o n . D i a g o n a l F l y  �  �        & e n t i t y . c r e a t u r e . m o b . c o m m o n . D i a g o n a l F l y   �  �        & e n t i t y . c r e a t u r e . m o b . c o m m o n . D i a g o n a l F l y   �  �        & e n t i t y . c r e a t u r e . m o b . c o m m o n . D i a g o n a l F l y   �  �        & e n t i t y . c r e a t u r e . m o b . c o m m o n . D i a g o n a l F l y   �  �        & e n t i t y . c r e a t u r e . m o b . c o m m o n . D i a g o n a l F l y   �  6        & e n t i t y . c r e a t u r e . m o b . c o m m o n . D i a g o n a l F l y   �  �        & e n t i t y . c r e a t u r e . m o b . c o m m o n . D i a g o n a l F l y   �  �        & e n t i t y . c r e a t u r e . m o b . c o m m o n . D i a g o n a l F l y   �          & e n t i t y . c r e a t u r e . m o b . c o m m o n . D i a g o n a l F l y   �  �        & e n t i t y . c r e a t u r e . m o b . c o m m o n . D i a g o n a l F l y   J           e n t i t y . i t e m . I t e m H o l d e r   �  �O o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . c o n s u m a b l e . s c r o l l . S c r o l l O f U p g r a d e        e n t i t y . i t e m . I t e m H o l d e r   �  �< o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . e n t i t i e s . C o i n        e n t i t y . c r e a t u r e . f x . H e a r t F x  �  U e n t i t y . c r e a t u r e . f x . H e a r t F x  �  0