   I   U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               	  	                                                                                                                                                                                                                                                                                    	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          	                                                                                                                                                                                                                                                          	                                                                                                                                                                                                                                                                  	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            	  	  	                                                                                                                                                          �   �  �  �   �  �  �                                                        	  	  	  	                                                                                                                                                        �   �   �   �   �   �   �                                                      	    	                                                                                                                         	  	  	    	                     �   �  �   �  �   �   �                                                     	    	                                                                                                                         	    	                     �  �   �  �  �   �   �                                                       	  	  	                                                                                                                                                        �   �   �   �   �  �   �                                                         	  	                                                                                                                                                          �  �   �  �   �  �   �                                                         	  	                                                                                                                                                           �   �   �   �   �   �   �                                                       	  	  	                                                                                                                                                          �   �   �  �  �   �   �                                                             	  	                                                                                                                                                                                                                                                                                                                                                                                                                                   	  	                                                                                                                                                                                                                                 	  	                                                                                                                                                                                                                                   	  	  	                                                                                                                                                                                                                             	                                                                                                    	                                                                                                                           	  	                                                                                                                                                                                                                        	  	                                                                                                                                                                                                                                                             	                                                                                                                                                                                                                               	  	                                                                                                                                                                                                                                               	  	  	  	                                                                                                                                                                                                                                              	  	  	  	                                                                                                                                                                                                                                               	    	  	                                                                                                                                                                                                                                                                          	                                                                                                                                                                                                                                                                 	  	                                                                      �  �  �   �   �   �   �  �   �                                                                                                                                                                                                                                   �   �   �   �   �   �   �  �   �                                                                                                                                                                                                                                 �   �   �   �  �   �   �   �   �                                                                                                                                                                                                                                      �   �   �   �   �   �  �  �   �                                                                                                                                                                                                                            �   �   �   �   �  �  �  �   �                                                                                                                                                                                                                                   �   �   �  �   �   �   �   �   �                                                                                                                                                                                                                                 �   �   �  �   �   �  �   �   �                                                                                                               	                                                                                                                 �  �  �  �   �   �  �   �  �                                                                                                                                                                                                                         �   �   �   �   �   �   �  �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   	           	                                                                                                                                                                                                                                       	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . S p i k e T r a p R o o m      2   #   C D o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . P a d R o o m            $ T o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . t r e a s u r e . C o r n e r l e s s T r e a s u r e R o o m      K   %   S N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . B o s s E n t r a n c e R o o m      /      8 R o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . V e r t i c a l S p i k e T r a p R o o m   6      G   # K o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . F i l l e d R o m b R o o m   3   :   ?   J H o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . b o s s . S i m p l e B o s s R o o m         "   / H o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s p e c i a l . N p c S a v e R o o m   ,      6    E o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . H e a r t R o o m            A o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . H a n d m a d e R o o m   #   =   3   F J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . H a l f R o o m C h a s m   &      1    P o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . t r e a s u r e . I s l a n d T r e a s u r e R o o m         &    N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . L i n e E n t r a n c e R o o m   #   -   ,   7  F o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s h o p . Q u a d S h o p R o o m   0   )   :   3S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . E m p t y C o n n e c t i o n R o o m      /      5 S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . E m p t y C o n n e c t i o n R o o m         &    S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . E m p t y C o n n e c t i o n R o o m   (      0   # M o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . R o l l i n g S p i k e R o o m   &   #   0   - O o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . C h a s m T u n n e l R o o m   0   #   8   ) J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . T u n n e l R o o m      C   #   K R o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . R i n g C o n n e c t i o n R o o m   '   	   ,    R o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . R i n g C o n n e c t i o n R o o m   ,      3       8                     	                                           	                                                         	       	      	      
      
      
      
      
         
                                                        
            
                                                      	                   
                              
   � e n t i t y . t r a p . R o l l i n g S p i k e  �  _��  �   ' e n t i t y . l e v e l . e n t i t i e s . c h e s t . W o o d e n C h e s t  �  � K o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . a c c e s s o r y . e q u i p p a b l e . F l i p p e r s        e n t i t y . l e v e l . e n t i t i e s . E x i t   �  8  e n t i t y . t r a p . R o l l i n g S p i k e    �    A�   e n t i t y . l e v e l . e n t i t i e s . D o o r     8   6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y A 1  e n t i t y . c r e a t u r e . n p c . T r a d e r     ` 
 
        d e n t i t y . c r e a t u r e . f x . H e a r t F x  C  � e n t i t y . c r e a t u r e . f x . H e a r t F x    �  e n t i t y . c r e a t u r e . f x . H e a r t F x  s  � e n t i t y . c r e a t u r e . f x . H e a r t F x  c  � e n t i t y . c r e a t u r e . f x . H e a r t F x  c  �' e n t i t y . l e v e l . e n t i t i e s . c h e s t . W o o d e n C h e s t       : o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . t o o l . M a t c h e s           e n t i t y . l e v e l . e n t i t i e s . E n t r a n c e  �    e n t i t y . l e v e l . e n t i t i e s . S l a b  !  � e n t i t y . i t e m . I t e m H o l d e r  "  �K o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . a c c e s s o r y . e q u i p p a b l e . R a g e R u n e       e n t i t y . l e v e l . e n t i t i e s . S l a b  �  � e n t i t y . i t e m . I t e m H o l d e r  �  �C o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . w e a p o n . s w o r d . C l a y m o r e         e n t i t y . l e v e l . e n t i t i e s . S l a b  !   e n t i t y . i t e m . I t e m H o l d e r     : o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . t o o l . M a t c h e s        e n t i t y . l e v e l . e n t i t i e s . S l a b  �   e n t i t y . i t e m . I t e m H o l d e r  �  I o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . w e a p o n . m a g i c . b o o k . C r a z y B o o k        e n t i t y . c r e a t u r e . n p c . S h o p k e e p e r  �  �          e n t i t y . t r a p . R o l l i n g S p i k e  �  _�   ��   e n t i t y . t r a p . R o l l i n g S p i k e  �  ��   A�   e n t i t y . t r a p . R o l l i n g S p i k e  �  _�   ��   e n t i t y . c r e a t u r e . f x . F i r e f l y  �   e n t i t y . c r e a t u r e . f x . F i r e f l y  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �    " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b   �  P" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b      0  e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y   �  A e n t i t y . c r e a t u r e . f x . F i r e f l y  Y  +" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  @  �  e n t i t y . c r e a t u r e . f x . F i r e f l y  G   ~ e n t i t y . c r e a t u r e . f x . F i r e f l y  �   � e n t i t y . c r e a t u r e . f x . F i r e f l y     ~" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b      P" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b      p  e n t i t y . c r e a t u r e . f x . F i r e f l y  c  o e n t i t y . c r e a t u r e . f x . F i r e f l y     � e n t i t y . c r e a t u r e . f x . F i r e f l y  B  � e n t i t y . c r e a t u r e . f x . F i r e f l y  Y  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  8" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b    �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  P  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  P  P " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  P  e n t i t y . c r e a t u r e . f x . F i r e f l y  �  ^" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  @ " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  P  @ e n t i t y . c r e a t u r e . f x . F i r e f l y  S   e n t i t y . c r e a t u r e . f x . F i r e f l y  �  Y e n t i t y . c r e a t u r e . f x . F i r e f l y  ]  1 e n t i t y . c r e a t u r e . f x . F i r e f l y  �  " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  [  � e n t i t y . c r e a t u r e . f x . F i r e f l y    v" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  P  ` e n t i t y . c r e a t u r e . f x . F i r e f l y  �   e n t i t y . c r e a t u r e . f x . F i r e f l y  �    e n t i t y . c r e a t u r e . f x . F i r e f l y  �  " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �     e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  \  k" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  p  @" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  p  � e n t i t y . c r e a t u r e . f x . F i r e f l y    `" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     p e n t i t y . c r e a t u r e . f x . F i r e f l y  �   � e n t i t y . c r e a t u r e . f x . F i r e f l y  �   � e n t i t y . c r e a t u r e . f x . F i r e f l y  �   � e n t i t y . c r e a t u r e . f x . F i r e f l y  	   � e n t i t y . c r e a t u r e . f x . F i r e f l y  �   � e n t i t y . c r e a t u r e . f x . F i r e f l y     � e n t i t y . l e v e l . e n t i t i e s . D o o r  �  @        4 e n t i t y . l e v e l . e n t i t i e s . D o o r  4       	  # A e n t i t y . l e v e l . e n t i t i e s . D o o r  4  0       # 3 e n t i t y . l e v e l . e n t i t i e s . D o o r    �         e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �         K e n t i t y . l e v e l . e n t i t i e s . D o o r    �         / e n t i t y . l e v e l . e n t i t i e s . D o o r  p  (        7 # e n t i t y . l e v e l . e n t i t i e s . D o o r  4        	  3 B e n t i t y . l e v e l . e n t i t i e s . D o o r  p  �         / e n t i t y . l e v e l . e n t i t i e s . D o o r    �        !  e n t i t y . l e v e l . e n t i t i e s . D o o r      �        2  e n t i t y . l e v e l . e n t i t i e s . D o o r  4  @    	   # D e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �     
   -  e n t i t y . l e v e l . e n t i t i e s . D o o r  �   �     
   *  e n t i t y . l e v e l . e n t i t i e s . D o o r  d       
   &  e n t i t y . l e v e l . e n t i t i e s . D o o r  d  �    
   &  e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �        ( - e n t i t y . l e v e l . e n t i t i e s . D o o r  �  (        , # e n t i t y . l e v e l . e n t i t i e s . D o o r    @       0 $ e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  �  �         e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  �  
      & e n t i t y . c r e a t u r e . m o b . h a l l . F r e e z i n g C l o w n  �  �         e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  �  
       e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �  y          e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f   �  �         # e n t i t y . c r e a t u r e . m o b . h a l l . I n v i s T h i e f   `  �          e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n   �  �         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f   �  �         % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t   �  �         e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t   w   
 
       e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n   P  p         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  0            # e n t i t y . c r e a t u r e . m o b . h a l l . I n v i s T h i e f    �          e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  �   �         e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t      � 
 
      % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  �           ' e n t i t y . c r e a t u r e . m o b . h a l l . S t a b b i n g K n i g h t     �        # e n t i t y . c r e a t u r e . m o b . h a l l . I n v i s T h i e f                e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  @           % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  %  �         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  p  p        # e n t i t y . c r e a t u r e . m o b . h a l l . I n v i s T h i e f  �  p         % e n t i t y . c r e a t u r e . m o b . h a l l . B u r n i n g C l o w n  P  @         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �  �          e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  H 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  `  p         # e n t i t y . c r e a t u r e . m o b . h a l l . I n v i s T h i e f  �  0          e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t      
 
      & e n t i t y . c r e a t u r e . m o b . h a l l . F r e e z i n g C l o w n     0        ' e n t i t y . c r e a t u r e . m o b . h a l l . S t a b b i n g K n i g h t  �  �         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  p  P         # e n t i t y . c r e a t u r e . m o b . h a l l . I n v i s T h i e f  �  P          e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �  p          e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  �  �         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  0            # e n t i t y . c r e a t u r e . m o b . h a l l . I n v i s T h i e f  0           # e n t i t y . c r e a t u r e . m o b . h a l l . I n v i s T h i e f  0            e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n      �        & e n t i t y . c r e a t u r e . m o b . h a l l . F r e e z i n g C l o w n              e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �  �         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �  p         % e n t i t y . c r e a t u r e . m o b . h a l l . B u r n i n g C l o w n  �  �         e n t i t y . i t e m . I t e m H o l d e r  �  �O o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . c o n s u m a b l e . s c r o l l . S c r o l l O f U p g r a d e        e n t i t y . i t e m . I t e m H o l d e r  �  �< o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . e n t i t i e s . C o i n        e n t i t y . i t e m . I t e m H o l d e r  �  �< o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . e n t i t i e s . C o i n        e n t i t y . i t e m . I t e m H o l d e r  p  \6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y B       