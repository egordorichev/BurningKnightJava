 S .         t                                                           J�        �        �        �        �       �       �                                                                   A�        �       �       �        �       �        �                �        �        �        �        �       �       �                A�        �       �       �        �       �        �                �        �        �        �       �       �       �                A�        �        �        �        �        �        �                 �        �        �        �        �        �        �                 A�        �        �       �        �        �        �                         �        �       �        �        �       �       �                A�       �       �        �        �       �       �                         �        �       �        �        �       �       �                 A�        �        �        �        �        �       �                �        �        �       �        �       �        �                A�        �        �       �        �       �       �                �       �        �        �        �        �        �                         ?        �        �        �        �       �        �       �                         �        �        �        �        �        �        �                =                                                                                                                                                      %                                                                                                                                                                                                                                                                            #                                                                                                                                                                                                                                                                                                                                                                 !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             (                                                                                                                                                                                                                                                                                                                   .                                                                                                                                                                                                                                                                          /                                                                                                                                                                                                                                 /                                                                                                                                                                                                                                                             /                                                                                                                                                                                                                                                                       /                                                                                                                                                                                                                                                     .                                                                                                                                                                                                                                                                   .                                                                                                                                                                                                                                                                  0                                  	                                                                    �D o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . B o m b R o o m   ' H o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . b o s s . S i m p l e B o s s R o o m      N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . B o s s E n t r a n c e R o o m M  Q  K o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . M i x e d S e c r e t R o o m )  1 N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . S m a l l A d d i t i o n R o o m   1  L o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . L i n e C i r c l e R o o m E  M   M o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . R o l l i n g S p i k e R o o m 1  E " M o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . C e n t e r S t r u c t R o o m   + , Q o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . t r e a s u r e . C o l l u m n T r e a s u r e R o o m     , P o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . S p i k e d T u n n e l R o o m     O o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . C h a s m T u n n e l R o o m +  1 # S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . E m p t y C o n n e c t i o n R o o m     (  		 

		

   I e n t i t y . i t e m . I t e m H o l d e r  3   `2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . i t e m . I t e m H o l d e r  3   `2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . i t e m . I t e m H o l d e r  3   `2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . l e v e l . e n t i t i e s . P o r t a l  �    e n t i t y . i t e m . I t e m H o l d e r  �   02 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . i t e m . I t e m H o l d e r  �   P6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C        e n t i t y . i t e m . I t e m H o l d e r  �   �6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C        e n t i t y . i t e m . I t e m H o l d e r  �   P2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . c r e a t u r e . f x . H e a r t F x  �   �% e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  �   0        % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  �   �         e n t i t y . l e v e l . e n t i t i e s . E n t r a n c e  �    e n t i t y . t r a p . R o l l i n g S p i k e  0  t    A�   e n t i t y . t r a p . R o l l i n g S p i k e  P  �    ��   e n t i t y . t r a p . R o l l i n g S p i k e  p  t    A�   e n t i t y . t r a p . R o l l i n g S p i k e  �  �    ��   e n t i t y . t r a p . R o l l i n g S p i k e  �  t    A�   e n t i t y . t r a p . R o l l i n g S p i k e  �  �    ��   e n t i t y . t r a p . R o l l i n g S p i k e  �  t    A�   e n t i t y . t r a p . R o l l i n g S p i k e    �    ��   e n t i t y . t r a p . R o l l i n g S p i k e  0  t    A�  ' e n t i t y . l e v e l . e n t i t i e s . c h e s t . W o o d e n C h e s t   �  ` K o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . a c c e s s o r y . e q u i p p a b l e . I c e B o o t s       " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b       �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  @   �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b      �  e n t i t y . c r e a t u r e . f x . F i r e f l y  �  '" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     0 e n t i t y . c r e a t u r e . f x . F i r e f l y  h   e n t i t y . c r e a t u r e . f x . F i r e f l y  �   � e n t i t y . c r e a t u r e . f x . F i r e f l y  �   �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b      �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  P  ` " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `   � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  @  @" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b      " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  @  " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  s  ;" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `   � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  9  Q" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  @  " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  @  0" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     @" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     `" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  @  p  e n t i t y . l e v e l . e n t i t i e s . D o o r  T  P       e n t i t y . l e v e l . e n t i t i e s . D o o r  �    < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . B u r n i n g K e y M  e n t i t y . l e v e l . e n t i t i e s . D o o r  �  P       e n t i t y . l e v e l . e n t i t i e s . D o o r    `     1  e n t i t y . l e v e l . e n t i t i e s . D o o r  T  @     E  e n t i t y . l e v e l . e n t i t i e s . D o o r    �     1  e n t i t y . l e v e l . e n t i t i e s . D o o r  T        ! e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �     +  e n t i t y . l e v e l . e n t i t i e s . D o o r   �  `      & e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �  @ 
 
        e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n     0        % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  �   �         e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �    
 
       e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �  � 
 
        e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  `  � 
 
        e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  �  P         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �  � 
 
        e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  �  P         e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n     �         e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  p    
 
        e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  `   
 
       e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  �  �         e n t i t y . c r e a t u r e . m o b . h a l l . C l o w n  �           e n t i t y . i t e m . I t e m H o l d e r  �  �< o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . e n t i t i e s . C o i n       