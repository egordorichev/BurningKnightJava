     !                                                                 	  	  	  	  	  	  	  	                    	  	  	  	  	  	  	  	  	              	  	  	  	  	  	  	  	                    	  	  	  	  	  	  	  	  	             	  	                                         	  	  	  	  	  	  	  	             	  	                                         	  	  	  	  	  	  	  	              	  	                                         	  	  	  	  	  	  	  	              	  	  	  	  	  	  	  	  	                  	  	  	  	  	  	  	  	  	              	  	  	  	  	  	  	  	  	                  	  	  	  	  	  	  	  	  	               	  	  	  	                            	  	  	  	  	  	  	  	  	              	  	  	                              	  	  	  	  	  	  	  	  	              	  	  	           	  	  	                  	  	  	  	  	  	  	  	  	               	  	  	          	  	  	                  	  	  	  	  	  	  	  	  	                             	  	                          	  	  	  	  	  	                                                                                                                                                                                                                                                                                                                                                              	                                                                     	               	                                                                      	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                8A o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . H a n d m a d e R o o m          e n t i t y . l e v e l . e n t i t i e s . E x i t   `   � # e n t i t y . l e v e l . e n t i t i e s . C l a s s S e l e c t o r   V   T@ o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . w e a p o n . s w o r d . S w o r d          w a r r i o r# e n t i t y . l e v e l . e n t i t i e s . C l a s s S e l e c t o r   �   VK o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . w e a p o n . m a g i c . M a g i c M i s s i l e W a n d          w i z a r d# e n t i t y . l e v e l . e n t i t i e s . C l a s s S e l e c t o r   q   QA o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . w e a p o n . g u n . R e v o l v e r            d    r a n g e r e n t i t y . c r e a t u r e . f x . F i r e f l y   �   ` e n t i t y . c r e a t u r e . f x . F i r e f l y  d  Q e n t i t y . c r e a t u r e . f x . F i r e f l y   X   � e n t i t y . c r e a t u r e . f x . F i r e f l y  I   ]" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b      �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b   �  p" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  p  p" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �