           \                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             
                                                                                                                                                                                                     	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              	                                              e< o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m     < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m  	   < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m    	 < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m  	   < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m     < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m  	   < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . S u b R o o m    	     O e n t i t y . l e v e l . e n t i t i e s . D o o r   �   �       e n t i t y . l e v e l . e n t i t i e s . D o o r   �          e n t i t y . l e v e l . e n t i t i e s . D o o r   �   �       	 e n t i t y . l e v e l . e n t i t i e s . E x i t      �  e n t i t y . l e v e l . e n t i t i e s . D o o r  D   �       e n t i t y . l e v e l . e n t i t i e s . D o o r  D          e n t i t y . l e v e l . e n t i t i e s . D o o r  `   �       	 e n t i t y . c r e a t u r e . n p c . U p g r a d e  `   � a f i r e _ f l o w e r e n t i t y . c r e a t u r e . n p c . U p g r a d e   @   � d	 w a l l _ b o o k e n t i t y . c r e a t u r e . n p c . U p g r a d e   P   � d t r i p l e _ b o o k e n t i t y . c r e a t u r e . n p c . U p g r a d e   `   � d c o n f e t t i _ g u n e n t i t y . c r e a t u r e . n p c . U p g r a d e   p   � d s h o v e l e n t i t y . c r e a t u r e . n p c . U p g r a d e   �   � d a i m _ b o o k e n t i t y . c r e a t u r e . n p c . U p g r a d e   �   � d c o n f e t t i _ g r e n a d e e n t i t y . c r e a t u r e . n p c . U p g r a d e   �   � d
 m a n a _ k n i f e e n t i t y . c r e a t u r e . n p c . U p g r a d e   �   P b s t a r t _ w i t h _ h e a l t h _ p o t i o n e n t i t y . c r e a t u r e . n p c . U p g r a d e   �   P b t o t a l l y _ s h o p e n t i t y . c r e a t u r e . n p c . U p g r a d e   �   D b e x t r a _ h e a r t e n t i t y . c r e a t u r e . n p c . U p g r a d e   P    c a p p l e e n t i t y . c r e a t u r e . n p c . U p g r a d e  �   � h	 d u n c e _ h a t e n t i t y . c r e a t u r e . n p c . U p g r a d e  �   � h m o a i _ h a t e n t i t y . c r e a t u r e . n p c . U p g r a d e  p   � h	 s k u l l _ h a t e n t i t y . c r e a t u r e . n p c . U p g r a d e  `   � h	 f u n g i _ h a t e n t i t y . c r e a t u r e . n p c . T r a d e r   o   � 
 
        c e n t i t y . c r e a t u r e . n p c . T r a d e r  `   � 
 
        h e n t i t y . c r e a t u r e . n p c . T r a d e r  Y   
 
        a e n t i t y . c r e a t u r e . n p c . T r a d e r   �   l 
 
       b e n t i t y . c r e a t u r e . n p c . T r a d e r   p   � 
 
        d e n t i t y . c r e a t u r e . n p c . U p g r a d e   �   D b b e t t e r _ c h e s t _ c h a n c e# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p   �   ~ s h o p - m a n i k e n# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p   �   � s h o p - t a r g e t# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p   �   z s h o p - s h i e l d s# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p  Q   � s h o p - c a r p e t# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p  �   �
 s h o p - s t a n d# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p  R   �
 s h o p - s t a n d# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p  �   �
 s h o p - s t a n d# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p  S   �
 s h o p - s t a n d( e n t i t y . l e v e l . e n t i t i e s . s h o p . S o l i d S h o p P r o p  k   �
 s h o p - s h e l f# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p   r  F	 s h o p - f r o g# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p   �  B s h o p - b a t# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p   d  C	 s h o p - b o n e# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p   �  B
 s h o p - s k u l l( e n t i t y . l e v e l . e n t i t i e s . s h o p . S o l i d S h o p P r o p   b  7
 s h o p - t a b l e( e n t i t y . l e v e l . e n t i t i e s . s h o p . S o l i d S h o p P r o p  r   s h o p - t a b l e _ 2 e n t i t y . c r e a t u r e . n p c . U p g r a d e  �   � a o b s i d i a n _ b o o t s e n t i t y . c r e a t u r e . n p c . U p g r a d e  p   � a c a m p f i r e _ i n _ a _ b o t t l e e n t i t y . c r e a t u r e . n p c . U p g r a d e  �   � a a n t i d o t e e n t i t y . c r e a t u r e . n p c . U p g r a d e   l    c b r e a d e n t i t y . c r e a t u r e . n p c . U p g r a d e   �    c m a p _ g r e e n p r i n t s e n t i t y . c r e a t u r e . n p c . U p g r a d e   �    c m a g i c _ m u s h r o o m# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p   .   �
 s h o p - b l o o d# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p   @   � s h o p - f r a m e _ b# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p   �   � s h o p - f r a m e _ b# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p   �   � s h o p - f r a m e _ a# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p   _   � s h o p - f r a m e _ a! e n t i t y . l e v e l . e n t i t i e s . H a t S e l e c t o r      h  ! e n t i t y . l e v e l . e n t i t i e s . H a t S e l e c t o r  @   h  ! e n t i t y . l e v e l . e n t i t i e s . H a t S e l e c t o r  `   h  ! e n t i t y . l e v e l . e n t i t i e s . H a t S e l e c t o r  �   h  ! e n t i t y . l e v e l . e n t i t i e s . H a t S e l e c t o r  `   H  ! e n t i t y . l e v e l . e n t i t i e s . H a t S e l e c t o r  �   I  ! e n t i t y . l e v e l . e n t i t i e s . H a t S e l e c t o r  @   H  ! e n t i t y . l e v e l . e n t i t i e s . H a t S e l e c t o r      H  # e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p  (   Q s h o p - c a r p e t# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p  �   ;
 s h o p - s t a n d# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p  �   {
 s h o p - s t a n d# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p     z
 s h o p - s t a n d# e n t i t y . l e v e l . e n t i t i e s . s h o p . S h o p P r o p     :
 s h o p - s t a n d e n t i t y . l e v e l . e n t i t i e s . B l o c k e r    ! e n t i t y . l e v e l . e n t i t i e s . H a t S e l e c t o r  0   X  ! e n t i t y . l e v e l . e n t i t i e s . H a t S e l e c t o r  P   X  ! e n t i t y . l e v e l . e n t i t i e s . H a t S e l e c t o r  p   X  ! e n t i t y . l e v e l . e n t i t i e s . H a t S e l e c t o r  0   q  ! e n t i t y . l e v e l . e n t i t i e s . H a t S e l e c t o r  p   r   e n t i t y . c r e a t u r e . f x . F i r e f l y  g   s e n t i t y . c r e a t u r e . f x . F i r e f l y  �   � e n t i t y . c r e a t u r e . f x . F i r e f l y  ~   � e n t i t y . c r e a t u r e . f x . F i r e f l y  �   � e n t i t y . c r e a t u r e . f x . F i r e f l y  f  	