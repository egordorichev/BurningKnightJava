    e n t i t y . c r e a t u r e . p l a y e r . P l a y e r   �   �        @ o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . w e a p o n . s w o r d . S w o r d                                A�         