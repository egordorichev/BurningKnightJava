 B y         \                                                                                                                                               *                                                                                                                                                                             )                                                                                                                                                                           )                                                                                                                                                                           )                                                                                                                                                                             )                                                                                                                                                                                )                                                                                                                                                                                 )                                                                                                                                                                                )                                                                                                                                                                                                                                                                                                                                                                                                             �       �       �       �        �       �        �                                                                                                                                                                                                 �        �        �       �        �       �        �                                                                                                                                                                                                                   �       �        �       �        �       �        �                                                                                                                                                                                                                                             �       �        �        �       �        �        �                                                                                                                                                                                                                         
                    �        �        �       �        �       �       �                                                                                                                                                                                                                                            �       �        �        �        �        �        �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      !                                                                                                                                                                                                                                      !                                                                                                                                                                                                                                     !                                                                                                                                                                                                                                   !                                                                                                                                                                                                                                   !                                                                                                                                                                                                                                !                                                                                                                                                                   5                                                                            7                                                                               7                                                                               7                                                                                +                 
                                                                               +                                                                                                                                                                     +                                                                                                                                                                  +                                                                                                                                                                +                                                                                                                                                                     +                                                                                                                                                                      +                                                                                                                                                                      +                                                                                                                                                                   +                                                                                                                                                                     +                                                                                                                                                                    +                                                                                                                                                                     +                                                                                                                                                                    +                                                                                                                                               7                                                                            7                                                                            7                                                                             7                                                                             7                                                                              6                                              3                                                            :                                                            :                                                            :                                                               5                                                                                                    4                                                                                                  4                                                                                              4                                                                                                       4                                                                                                        4                                                                                                       4                                                                                                  4                                                                                              4                                                                                                4                                                                                               4                                                                                              4                                                                                             4                                                                                                  4                                                                                                   4                                                                                                      4                                                                                          5                      �        �        �        �       �       �        �        �        �                 5                       �        �        �        �       �       �       �        �        �                         1                                      �        �        �        �       �       �        �       �        �                 0                                                    �        �        �        �        �       �        �        �        �                         "                                 	                                            �        �        �        �        �        �        �        �        �                        "                                  	                                                        �        �        �       �       �        �        �        �       �                        )                                                                                                                        $                                                                                                ,                                                                                            "                                                                                                                                                                                                  !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ,                                                                                                                                                              -                                                                                                                                                                          +                                                                                                                                                                                       ,                                                                                                                                                                       ,                                                                                                                                                                           -                                                                                                                                                                 -                                                                                                                                                                 ,                                                                                                                                                                        -                                                                                                                                                                   -                                                                                                                                                                   -                                                                                                                                                                      ,                                                                                                                                                             -                                                                                                                                                             ,                                                                                                                                                                              +                                                                                                                              �K o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . i t e m . B r o k e L i n e I t e m R o o m ( 2 4 B H o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . F l o o d e d R o o m  L - a T o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . t r e a s u r e . C o r n e r l e s s T r e a s u r e R o o m #  / ( J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . G o l d S e c r e t R o o m + B 5 IH o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . b o s s . S i m p l e B o s s R o o m  a ) w L o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . L i n e C i r c l e R o o m 2  :   D o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . P a d R o o m   2  J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . C a v y C h a s m R o o m /  8 . N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . B o s s E n t r a n c e R o o m 4  8  G o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . G a r d e n R o o m  L  a I o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s h o p . C l a s s i c S h o p R o o m  a  h K o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . M i x e d S e c r e t R o o m 8 	 @ S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . C h a s m C o n n e c t i o n R o o m + . 1 2 J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . T u n n e l R o o m ) B + E J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . T u n n e l R o o m $ E + L J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . T u n n e l R o o m  F  L *   	 			
		
	  	   O e n t i t y . l e v e l . e n t i t i e s . S l a b  �  �' e n t i t y . l e v e l . e n t i t i e s . c h e s t . W o o d e n C h e s t  �    B o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . w e a p o n . s w o r d . B u t c h e r          e n t i t y . i t e m . I t e m H o l d e r  �  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r    �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  3  P2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �  P2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  C  P2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d       % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t    p        % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  0  `         e n t i t y . l e v e l . e n t i t i e s . E n t r a n c e  a  :  e n t i t y . l e v e l . e n t i t i e s . E x i t  `   �  e n t i t y . l e v e l . e n t i t i e s . S l a b   2  8 e n t i t y . i t e m . I t e m H o l d e r   4  ?2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b       e n t i t y . l e v e l . e n t i t i e s . S l a b   R  8 e n t i t y . i t e m . I t e m H o l d e r   T  ?6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C       e n t i t y . l e v e l . e n t i t i e s . S l a b   r  8 e n t i t y . i t e m . I t e m H o l d e r   u  N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . a c c e s s o r y . e q u i p p a b l e . V a m p i r e R i n g       e n t i t y . l e v e l . e n t i t i e s . S l a b   �  8 e n t i t y . i t e m . I t e m H o l d e r   �  : o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . I n f i n i t e B o m b       e n t i t y . l e v e l . e n t i t i e s . S l a b   �  8 e n t i t y . i t e m . I t e m H o l d e r   �  >F o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . p e t . o r b i t a l . J e l l y O r b i t a l       e n t i t y . l e v e l . e n t i t i e s . S l a b   �  8 e n t i t y . i t e m . I t e m H o l d e r   �  AJ o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . a c c e s s o r y . e q u i p p a b l e . T e c h E y e      $ e n t i t y . c r e a t u r e . n p c . O r a n g e S h o p k e e p e r   @             e n t i t y . i t e m . I t e m H o l d e r   �  !2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �   �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . i t e m . I t e m H o l d e r  �   �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . i t e m . I t e m H o l d e r  �   �6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C        e n t i t y . i t e m . I t e m H o l d e r  �   �6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C        e n t i t y . i t e m . I t e m H o l d e r  �   �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �   �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . c r e a t u r e . f x . H e a r t F x  �   � e n t i t y . c r e a t u r e . f x . F i r e f l y  #  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  0   e n t i t y . c r e a t u r e . f x . F i r e f l y  2  f" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �    e n t i t y . c r e a t u r e . f x . F i r e f l y  �  C e n t i t y . c r e a t u r e . f x . F i r e f l y  C   " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  `" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b       e n t i t y . c r e a t u r e . f x . F i r e f l y  #  � e n t i t y . c r e a t u r e . f x . F i r e f l y  ]  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     � " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  p  � e n t i t y . c r e a t u r e . f x . F i r e f l y  j   � e n t i t y . c r e a t u r e . f x . F i r e f l y  Q  � e n t i t y . c r e a t u r e . f x . F i r e f l y  k  j" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �   " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b      e n t i t y . c r e a t u r e . f x . F i r e f l y  �  @" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  @" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  P  �  e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . l e v e l . e n t i t i e s . D o o r  �       * B e n t i t y . l e v e l . e n t i t i e s . D o o r  �       / 2 e n t i t y . l e v e l . e n t i t i e s . D o o r  P  �     % L e n t i t y . l e v e l . e n t i t i e s . D o o r  0       # a e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �      L e n t i t y . l e v e l . e n t i t i e s . D o o r  �  @     T e n t i t y . l e v e l . e n t i t i e s . D o o r  �  0    / # e n t i t y . l e v e l . e n t i t i e s . D o o r  `   �   < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . B u r n i n g K e y 6  e n t i t y . l e v e l . e n t i t i e s . D o o r  $  `    2  e n t i t y . l e v e l . e n t i t i e s . D o o r  @  h     4  e n t i t y . l e v e l . e n t i t i e s . D o o r     h     0  e n t i t y . l e v e l . e n t i t i e s . D o o r     �     0 . e n t i t y . l e v e l . e n t i t i e s . D o o r   �     6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C  a e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �      L% e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t   �  �         e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  ]  � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  O  s  
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  <  �  
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  i  s 
 
       e n t i t y . i t e m . I t e m H o l d e r  n   �< o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . e n t i t i e s . C o i n        e n t i t y . i t e m . I t e m H o l d e r  �   $B o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . p l a n t . s e e d . G r a s s S e e d        e n t i t y . c r e a t u r e . f x . H e a r t F x     � e n t i t y . i t e m . I t e m H o l d e r    �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d       