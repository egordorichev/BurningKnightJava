 ` �    �                          X                                                             P                                                                  P                                	                         P                                	   	   	      	                Q                                   	   	                    Q                                                             Q                                                             Q                                                             P                                                                             N                                                                                 M                                                                        M                                                                             &         &                                                                         #                                                                                                                       !                                                                                                                               #                                                                                                                                                    #                                                                                                                                                       #                                                                                                                                                                #                                                                                                                                                                        #                                                                                                                                                                                            "                                                                                                                                                                "                                                                                                                                         "                                                                                                                                                                                     #                                                                                                                                                                                                              ,                                                                                                                                                                               .                                                                                                                                                               .                                                                                                                                             4                                                                                                                                                          5                                                                                                                                           5                                                                                                                                                   5                                                                                                                     :                                                                                                                                                   3                                                                                                                                                        6                                                                                                                          H                                                    L                                                                                         I                                                                                           I                                                                                           I                                                                  L                                   L                                                                     J                                                K                                                                  H         	                                           K                                                                 P                                                   I                                                                  G                                            J                                          	   	        M                                            	   	                    H                                             	   	   	                    H                                                                                                H                                                                                             H                                                                                          I                                  W                         �    �   �    �    �   �   �    �         Q              �    �    �    �    �   �    �    �            P              �   �                 �   �         B                                           �    �         �    �         �   �         C                                                                             �    �        �    �        �    �         C                                                                         �    �                  �    �         B                                                   �   �    �    �    �    �    �   �         B                                                          �    �   �    �    �    �   �   �             A                                                                                                B                     	                 	            R                                         	        R                                                       P                                       	                 Q                                       Z                         Y                             Y                                 X                                 X                             Y                                 R                                                6                                                                                                                               ;                                                                                                                        ;                                                                                             ;                                                                                                                                            ;                                                                                                                              :                                                                                                                                                   ;                                                                                                                                     ;                                                                                                                                                :                                                                                                                                                9                                                                                                                                                   ;                                                                                                        :                                                                                 H                                                                                      G                                                                                                   H                                                                                     H                                                                                                    C                                                                        A                                   	                                                             A                                                                                          F                                                                                      F                                                                                                       F                                                                                                     F                                                                                                         F                                                                                                         F                                                                                                          G                                                                                                  D                                                                                                                     F                                                                                                       @                                                                                          C                                                                             E                                                                                      B                                                                                        A                                                                                         B                                                                                              A                                                                          C                                                                 J                                                                 J                                                                      I                                                                   D                                                            C                                                                                                      C                                                                                                   C                                                                                           G                                                                       N                                                      N                                                                                     L                                                                           U                                                                  O                                                                             M                                                                         N                                                                             M                                                                       N                                     	                               N                         	      	                                 N                             	                                       M                                                                   N                                                                     N                                                                         M                                                                    N                                                                     N                                                                    N                                                                           M                                                                        N                                                                       M                                                                          N                                                                         M                                            	   	                            M                                                                            N                                               6N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . M i s s i n g C o r n e r R o o m D ! R * H o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . C o l l u m n R o o m '  > ) K o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . S i d e C h a s m s R o o m E  T  J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . E n t r a n c e R o o m  r  {  N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . B o s s E n t r a n c e R o o m  {  � K o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . F i l l e d R o m b R o o m  d $ r N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . t r e a s u r e . M a z e T r e a s u r e R o o m  T $ d R o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . V e r t i c a l S p i k e T r a p R o o m 9 * P > H o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s p e c i a l . N p c S a v e R o o m  r $ ~ H o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . b o s s . S i m p l e B o s s R o o m F  X ! G o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . C i r c l e R o o m  � ( � D o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . P a d R o o m , S 9 ^ S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . t r e a s u r e . B r o k e L i n e T r e a s u r e R o o m   '   K o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . i t e m . B r o k e L i n e I t e m R o o m 0 B > L J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . G o l d S e c r e t R o o m D > M GS o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . E m p t y C o n n e c t i o n R o o m $ ^ , f R o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . R i n g C o n n e c t i o n R o o m ' W , ^ O o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . C h a s m T u n n e l R o o m 6 L < S R o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . R i n g C o n n e c t i o n R o o m > > D D O o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . C h a s m T u n n e l R o o m >  F  S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . E m p t y C o n n e c t i o n R o o m 7  >  J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . T u n n e l R o o m  {  � S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . C h a s m C o n n e c t i o n R o o m $ f ( n S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . C h a s m C o n n e c t i o n R o o m $ n , v <  		 
	 		

	
   � e n t i t y . l e v e l . e n t i t i e s . E n t r a n c e  !  j  e n t i t y . l e v e l . e n t i t i e s . E x i t   �  � ! e n t i t y . l e v e l . e n t i t i e s . c h e s t . M i m i c  �  �           e n t i t y . t r a p . R o l l i n g S p i k e  �  �    A�   e n t i t y . l e v e l . e n t i t i e s . D o o r  �  H   6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y A  u e n t i t y . c r e a t u r e . n p c . T r a d e r  �  � 
 
        d! e n t i t y . l e v e l . e n t i t i e s . c h e s t . M i m i c    �          e n t i t y . l e v e l . e n t i t i e s . S l a b  p  p e n t i t y . i t e m . I t e m H o l d e r  r  rO o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . c o n s u m a b l e . s c r o l l . S c r o l l O f U p g r a d e        e n t i t y . i t e m . I t e m H o l d e r  �   2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �  2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �  @2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �  `2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d       " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  P   " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �   � e n t i t y . c r e a t u r e . f x . F i r e f l y  �   � e n t i t y . c r e a t u r e . f x . F i r e f l y  !  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  P" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  p  `" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b    �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     � " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     � " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  @  �  e n t i t y . c r e a t u r e . f x . F i r e f l y  (  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  r" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  P" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  P  P " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  p" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b    � " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  0  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  0  � " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  0  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `   e n t i t y . c r e a t u r e . f x . F i r e f l y  �  0 e n t i t y . c r e a t u r e . f x . F i r e f l y  %  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     ` e n t i t y . c r e a t u r e . f x . F i r e f l y  C  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  p    " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  p    e n t i t y . c r e a t u r e . f x . F i r e f l y  �  	n e n t i t y . c r e a t u r e . f x . F i r e f l y    	 e n t i t y . c r e a t u r e . f x . F i r e f l y  �  	@ e n t i t y . c r e a t u r e . f x . F i r e f l y  �  {" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  p  @ e n t i t y . c r e a t u r e . f x . F i r e f l y  -  � e n t i t y . c r e a t u r e . f x . F i r e f l y  <  g e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  ;  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  @  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  @  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  r e n t i t y . c r e a t u r e . f x . F i r e f l y  u  C e n t i t y . c r e a t u r e . f x . F i r e f l y  v  	 e n t i t y . c r e a t u r e . f x . F i r e f l y  |  ] e n t i t y . c r e a t u r e . f x . F i r e f l y  z  '" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  P  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  P e n t i t y . c r e a t u r e . f x . F i r e f l y  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �   e n t i t y . c r e a t u r e . f x . F i r e f l y  8  � e n t i t y . c r e a t u r e . f x . F i r e f l y  ?  � e n t i t y . c r e a t u r e . f x . F i r e f l y  M  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  P  p e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  ?  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  p  p" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  p  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �   e n t i t y . l e v e l . e n t i t i e s . D o o r  p  �         G * e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �        8  e n t i t y . l e v e l . e n t i t i e s . D o o r  t  �       '  e n t i t y . l e v e l . e n t i t i e s . D o o r  �   �      	  M  e n t i t y . l e v e l . e n t i t i e s . D o o r     �   < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . B u r n i n g K e y  { e n t i t y . l e v e l . e n t i t i e s . D o o r     �         { e n t i t y . l e v e l . e n t i t i e s . D o o r  D  �       $ k e n t i t y . l e v e l . e n t i t i e s . D o o r  �  8         d e n t i t y . l e v e l . e n t i t i e s . D o o r     �        @ > e n t i t y . l e v e l . e n t i t i e s . D o o r  D  0       $ s e n t i t y . l e v e l . e n t i t i e s . D o o r  d  �    	   F  e n t i t y . l e v e l . e n t i t i e s . D o o r  p  (     
    � e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �       , ] e n t i t y . l e v e l . e n t i t i e s . D o o r  �  (        8 S e n t i t y . l e v e l . e n t i t i e s . D o o r  �  0       > C e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �        : L e n t i t y . l e v e l . e n t i t i e s . D o o r  p  �        ' n e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  @ 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  r  @ 
 
      % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  �  H         e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  `  P 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  ( 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  b 
 
      % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  `  �        e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �    
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �   � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �   � 
 
      e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �   � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t     � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t     � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t    � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  � 
 
      % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  �  �        % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t    �        % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  �  �         e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  ` 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  	P 
 
      % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t     p         e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t    � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  	4 
 
      % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t    O        % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  �  s        % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  d  z         e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  `  � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  c  � 
 
      % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  @  �        % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t  �  i         e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  q  M 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  �  p 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  y  x 
 
       e n t i t y . i t e m . I t e m H o l d e r   �  �< o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . e n t i t i e s . C o i n        e n t i t y . i t e m . I t e m H o l d e r  b  �6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y A       