    
 F i r e P o t i o n G R E E N  H e a l i n g P o t i o n Y E L L O W  I n v i s i b i l i t y P o t i o n B L U E  P o i s o n P o t i o n R E D  R e g e n e r a t i o n P o t i o n O R A N G E     B�      