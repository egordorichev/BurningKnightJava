 9 y         U                                  -                                                                                                    +                                                                                                      +                                                                                         +                                                                                                      +                                                                                                        +                                                                                                       +                                                                                                        +                                                                                                      +                                                            +                                                                                                +                                                                                                +                                                                                  0                                                                0                                                                                &                                                                                                            "                                                                                                          "                                                                                                                                              "                                                                                                                                                                      "                                                                                                                                                                !                                                                                                                        (                                                                                                                       (                                                                                                                     (                                                                                                                                                                                                           �       �        �       �        �        �       �       �       �                                                                                                                   �       �        �       �        �       �        �       �        �                                                                                                                                                                    �       �       �        �        �       �        �        �       �                                                                                                                                                                           �        �        �        �       �       �        �        �       �                                                                                                                                                                               �        �       �        �       �        �        �        �       �                                                                                                                                                                                �        �       �        �        �        �        �        �        �                                                                                                                                                                                          �        �        �        �       �       �       �       �        �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           !                                                                                                                                                                        !                                                                                                                                                                       !                                                                                                                                                                    !                                                                                                                                                                      !                                                                                          $                                                      2                                                      2                                                      2                                                     2                                       3                                                                         /                                                                          /                                                                         /                                                                          /                                                                         ,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   $                                                                                                                                                                                 "                                                                                                                                                                                 $                                                                                                                                                                       $                                                                                                                                                                     $                                                                                                                                                                   $                                                                                                                                                                            #                                                                                                                                                                     #                                                                                                                                                                             &                                                                                                                      %        �       �        �        �        �        �                                                                               $�        �        �        �        �        �                                                                         $        �       �        �        �        �       �                                                                                           �       �        �        �       �        �                                                                                                                                                  �        �        �        �        �       �                                                                                                                                                  �       �       �        �        �       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  !                                                                                                                                                                                         !                                                                                                                                                                                                 "                                                                                                                                                                                                 !                                                                                                                                                                                                 !                                                                                                                                                                                         !                                                                                                                                                                                                                                                                                                                                                                                                       !                                                                                                                                                                                               (                                                                                             �N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . M i s s i n g C o r n e r R o o m  4  E N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . B o s s E n t r a n c e R o o m 2  6  H o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . B i g H o l e R o o m   5 ( H o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . b o s s . S i m p l e B o s s R o o m  a % w I o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s h o p . C l a s s i c S h o p R o o m  H , O J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . R e c t F l o o r R o o m  E  Y P o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . t r e a s u r e . I s l a n d T r e a s u r e R o o m % c 1 m H o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s p e c i a l . N p c S a v e R o o m   (  J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . C a v y C h a s m R o o m  4 % G K o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . M i x e d S e c r e t R o o m  Y  `D o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . B o m b R o o m    !L o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . L i n e C i r c l e R o o m .  7   S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . E m p t y C o n n e c t i o n R o o m " ( ' - S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . E m p t y C o n n e c t i o n R o o m # - + 4 S o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . C h a s m C o n n e c t i o n R o o m  Y  a J o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . T u n n e l R o o m  G  L O o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . C h a s m T u n n e l R o o m % \ - c R o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . R i n g C o n n e c t i o n R o o m (  .  P o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . S p i k e d T u n n e l R o o m !  (  *  
 	 	
   Y e n t i t y . l e v e l . e n t i t i e s . P o r t a l  @    e n t i t y . l e v e l . e n t i t i e s . S l a b  �  � e n t i t y . i t e m . I t e m H o l d e r  �  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . l e v e l . e n t i t i e s . S l a b    � e n t i t y . i t e m . I t e m H o l d e r    �L o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . a c c e s s o r y . e q u i p p a b l e . O l d M a n u a l        e n t i t y . l e v e l . e n t i t i e s . S l a b  "  � e n t i t y . i t e m . I t e m H o l d e r  #  �B o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . c o n s u m a b l e . f o o d . P i l l        e n t i t y . l e v e l . e n t i t i e s . S l a b  B  � e n t i t y . i t e m . I t e m H o l d e r  C  �? o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . w e a p o n . g u n . P i s t o l             e n t i t y . l e v e l . e n t i t i e s . S l a b  b  � e n t i t y . l e v e l . e n t i t i e s . S l a b  �  � e n t i t y . l e v e l . e n t i t i e s . S l a b  �  �' e n t i t y . l e v e l . e n t i t i e s . c h e s t . W o o d e n C h e s t  �  � L o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . w e a p o n . t h r o w i n g . T h r o w i n g D a g g e r           e n t i t y . l e v e l . e n t i t i e s . D o o r      8   6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C "  e n t i t y . c r e a t u r e . n p c . T r a d e r      p 
 
        d e n t i t y . i t e m . I t e m H o l d e r   c  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . i t e m . I t e m H o l d e r   c  �6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C        e n t i t y . i t e m . I t e m H o l d e r   s  �6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C        e n t i t y . i t e m . I t e m H o l d e r   �  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . c r e a t u r e . f x . H e a r t F x   �  �  e n t i t y . c r e a t u r e . f x . H e a r t F x   �  �  e n t i t y . i t e m . I t e m H o l d e r  �  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . i t e m . I t e m H o l d e r  �  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . i t e m . I t e m H o l d e r  �  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . i t e m . I t e m H o l d e r  �  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . l e v e l . e n t i t i e s . E n t r a n c e  1  j  e n t i t y . c r e a t u r e . f x . F i r e f l y  J   e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y   �  � e n t i t y . c r e a t u r e . f x . F i r e f l y   f  | e n t i t y . c r e a t u r e . f x . F i r e f l y  '  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b      `" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b      � " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  P  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  `" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b      P" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b      � " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  @   � e n t i t y . c r e a t u r e . f x . F i r e f l y   q  � e n t i t y . c r e a t u r e . f x . F i r e f l y   w  � e n t i t y . c r e a t u r e . f x . F i r e f l y    � e n t i t y . c r e a t u r e . f x . F i r e f l y  <  � e n t i t y . c r e a t u r e . f x . F i r e f l y  E  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `  @ e n t i t y . c r e a t u r e . f x . F i r e f l y  \  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  p    e n t i t y . c r e a t u r e . f x . F i r e f l y  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  p  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  p  � " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �   e n t i t y . c r e a t u r e . f x . F i r e f l y  �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `     e n t i t y . c r e a t u r e . f x . F i r e f l y  k  / e n t i t y . c r e a t u r e . f x . F i r e f l y  _   e n t i t y . c r e a t u r e . f x . F i r e f l y  O  &" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  p   � e n t i t y . l e v e l . e n t i t i e s . D o o r   �  H       E e n t i t y . l e v e l . e n t i t i e s . D o o r  @  (   < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . B u r n i n g K e y 4  e n t i t y . l e v e l . e n t i t i e s . D o o r     �      0  e n t i t y . l e v e l . e n t i t i e s . D o o r  P  x      % ( e n t i t y . l e v e l . e n t i t i e s . D o o r  T        % b e n t i t y . l e v e l . e n t i t i e s . D o o r  P         a e n t i t y . l e v e l . e n t i t i e s . D o o r  �  �      I e n t i t y . l e v e l . e n t i t i e s . D o o r  d  `      F e n t i t y . l e v e l . e n t i t i e s . D o o r     �       Y e n t i t y . l e v e l . e n t i t i e s . D o o r  d  �      H e n t i t y . l e v e l . e n t i t i e s . D o o r  �  (      + c e n t i t y . l e v e l . e n t i t i e s . D o o r  `   �      &  e n t i t y . l e v e l . e n t i t i e s . D o o r  @  8      $ 4 e n t i t y . l e v e l . e n t i t i e s . D o o r  �  h       G e n t i t y . l e v e l . e n t i t i e s . D o o r  �  @     .  e n t i t y . l e v e l . e n t i t i e s . D o o r  �  @     (  e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f   �  p 
 
        e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t     � 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f   �    
 
        e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  P  � 
 
        e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t  P  0 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t   p    
 
       e n t i t y . c r e a t u r e . m o b . h a l l . K n i g h t    p 
 
       e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f   �  P 
 
       % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t   0  �        % e n t i t y . c r e a t u r e . m o b . h a l l . R a n g e d K n i g h t   �  �         e n t i t y . i t e m . I t e m H o l d e r   �  �O o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . c o n s u m a b l e . s c r o l l . S c r o l l O f U p g r a d e        e n t i t y . c r e a t u r e . f x . H e a r t F x    � 