   i         .                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �       �        �        �        �        �        �                                                                                               �        �       �        �       �       �        �                                                                                                    �        �        �       �        �        �        �                                                                                              �        �       �        �        �        �       �                                                                                                       �        �        �        �        �        �        �                                                                                                �        �        �       �        �        �       �                                                                                                       �        �       �       �        �        �        �                                                                                        �        �        �        �        �        �        �                                                                                                �        �        �        �        �        �        �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �        �        �       �        �        �       �        �       �                                                                                                               
�        �        �       �       �       �        �        �        �                                                                                                                        �        �       �       �        �       �       �        �        �                                                                                                                                       �        �       �        �       �       �        �       �        �                                                                                                                        �       �       �        �        �        �        �        �       �                                                                                                                         �       �       �        �        �        �        �       �        �                                                                                                                         	�        �        �        �        �        �        �        �        �                                                                                                                 	�        �       �        �        �        �        �        �       �                                                                                                                                   �        �        �        �       �       �       �        �        �                                                                                                                          	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    IJ o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . G o l d S e c r e t R o o m    &Q o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . t r e a s u r e . C o l l u m n T r e a s u r e R o o m  _  g H o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . b o s s . S i m p l e B o s s R o o m  /  E N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . B o s s E n t r a n c e R o o m     L o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . e n t r a n c e . L i n e C i r c l e R o o m      M o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . D o u b l e C o r n e r R o o m  K  _ D o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . P a d R o o m     N o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . r e g u l a r . S m a l l A d d i t i o n R o o m    / K o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . s e c r e t . M i x e d S e c r e t R o o m  R  \R o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . R i n g C o n n e c t i o n R o o m     P o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . S p i k e d T u n n e l R o o m  E  K R o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . l e v e l . r o o m s . c o n n e c t i o n . R i n g C o n n e c t i o n R o o m  _  e  

		 		

   A e n t i t y . i t e m . I t e m H o l d e r  �  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  �  2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . i t e m . I t e m H o l d e r  s  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d       ! e n t i t y . l e v e l . e n t i t i e s . c h e s t . M i m i c     0           e n t i t y . l e v e l . e n t i t i e s . P o r t a l      (  e n t i t y . l e v e l . e n t i t i e s . E n t r a n c e     �  e n t i t y . i t e m . I t e m H o l d e r   S  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . B o m b        e n t i t y . i t e m . I t e m H o l d e r   �  �6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C        e n t i t y . i t e m . I t e m H o l d e r   C  �6 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . K e y C        e n t i t y . i t e m . I t e m H o l d e r   c  �2 o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . G o l d        e n t i t y . c r e a t u r e . f x . H e a r t F x   #  � e n t i t y . c r e a t u r e . f x . F i r e f l y  �  5 e n t i t y . c r e a t u r e . f x . F i r e f l y  �  F e n t i t y . c r e a t u r e . f x . F i r e f l y  �  +" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b   �  `  e n t i t y . c r e a t u r e . f x . F i r e f l y   �  m" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b      " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     @ e n t i t y . c r e a t u r e . f x . F i r e f l y   �   t" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b   �   `" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  0   `" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  0   � e n t i t y . c r e a t u r e . f x . F i r e f l y  Z  x e n t i t y . c r e a t u r e . f x . F i r e f l y   �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  `  0" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b   �  p" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b     �  e n t i t y . c r e a t u r e . f x . F i r e f l y   �   �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b    " e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  �  � e n t i t y . c r e a t u r e . f x . F i r e f l y  <  � e n t i t y . c r e a t u r e . f x . F i r e f l y   �   e n t i t y . c r e a t u r e . f x . F i r e f l y  4  � e n t i t y . c r e a t u r e . f x . F i r e f l y   �  N e n t i t y . c r e a t u r e . f x . F i r e f l y  0  � e n t i t y . c r e a t u r e . f x . F i r e f l y  :  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b  @  � e n t i t y . c r e a t u r e . f x . F i r e f l y   �  � e n t i t y . c r e a t u r e . f x . F i r e f l y   �  �" e n t i t y . l e v e l . e n t i t i e s . d e c o r . C o b w e b   �  ` e n t i t y . c r e a t u r e . f x . F i r e f l y  �  > e n t i t y . l e v e l . e n t i t i e s . D o o r  d  @      d e n t i t y . l e v e l . e n t i t i e s . D o o r   �  H       E e n t i t y . l e v e l . e n t i t i e s . D o o r   �  �       / e n t i t y . l e v e l . e n t i t i e s . D o o r     H   < o r g . r e x c e l l e n t g a m e s . b u r n i n g k n i g h t . e n t i t y . i t e m . k e y . B u r n i n g K e y   e n t i t y . l e v e l . e n t i t i e s . D o o r   �   �        e n t i t y . l e v e l . e n t i t i e s . D o o r   �  �       K e n t i t y . l e v e l . e n t i t i e s . D o o r  p  �       _ e n t i t y . l e v e l . e n t i t i e s . D o o r  0  �        e n t i t y . l e v e l . e n t i t i e s . D o o r  @  �       ' e n t i t y . c r e a t u r e . m o b . d e s e r t . A r c h e o l o g i s t    P 
 
      ' e n t i t y . c r e a t u r e . m o b . d e s e r t . A r c h e o l o g i s t  @   
 
       e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  @    
 
        e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f   �  @ 
 
       ' e n t i t y . c r e a t u r e . m o b . d e s e r t . A r c h e o l o g i s t     � 
 
      # e n t i t y . c r e a t u r e . m o b . d e s e r t . S k e l e t o n   �  �       ' e n t i t y . c r e a t u r e . m o b . d e s e r t . A r c h e o l o g i s t    P 
 
        e n t i t y . c r e a t u r e . m o b . d e s e r t . M u m m y  p   
 
       e n t i t y . c r e a t u r e . m o b . h a l l . T h i e f  �    
 
       ' e n t i t y . c r e a t u r e . m o b . d e s e r t . A r c h e o l o g i s t  P  ` 
 
      ' e n t i t y . c r e a t u r e . m o b . d e s e r t . A r c h e o l o g i s t     ` 
 
        e n t i t y . c r e a t u r e . m o b . d e s e r t . M u m m y     � 
 
        e n t i t y . c r e a t u r e . m o b . d e s e r t . M u m m y   �   
 
     ' e n t i t y . c r e a t u r e . m o b . d e s e r t . A r c h e o l o g i s t    � 
 
        e n t i t y . c r e a t u r e . m o b . d e s e r t . M u m m y  @  � 
 
      