    s e t t i n g s _ g o r e t r u e n u m _ b u l l e t s _ r e f l e c t e d 5 s e t t i n g s _ q u a l i t y 1 U N L O C K _ B L A C K _ H E A R T t r u e h i d e _ m i n i m a p t r u e s e t t i n g s _ v s y n c t r u e
 l a s t _ c l a s s 0 s e t t i n g s _ u i s f x t r u e s e t t i n g s _ b l o o d t r u e s e t t i n g s _ f u l l s c r e e n f a l s e s e t t i n g s _ c u r s o r c u r s o r - s t a n d a r t s e t t i n g s _ r o t a t e _ c u r s o r t r u e U P G R A D E _ A C H I E V E M E N T t r u e s e t t i n g s _ s f x 0 . 7 5 s e t t i n g s _ m u s i c 0 . 5 E Q U I P _ A C C E S S O R Y _ A C H I E V E M E N T t r u e s e t t i n g s _ s c r e e n s h a k e 0 . 7 T U T O R I A L _ D O N E _ A C H I E V E M E N T t r u e